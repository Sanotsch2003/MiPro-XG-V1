    signal ram : ram_type :=(
        0 => "11111101110000000001001100000000",
        1 => "11111101111010000000000000001100",
        2 => "11111001000000000000110000000000",
        3 => "11111101110111100001000000000001",
        4 => "11111101111000000101111101001100",
        5 => "11111001000000000000110000010001",
        6 => "11110000100000000000000000000001",
        7 => "11111101110000000001010000000000",
        8 => "11111101111010000000000000001100",
        9 => "11111001000000000000110000000000",
        10 => "11111101110000000000000000100001",
        11 => "11110000100000000000000000000001",
        12 => "11111101110000000000101000000000",
        13 => "11111101111010000000000000001100",
        14 => "11111001000000000000110000000000",
        15 => "11111101110001001000010010000001",
        16 => "11111101111000000001111010001100",
        17 => "11111001000000000000110000010001",
        18 => "11110000100000000000000000000001",
        19 => "11111101110000000001010010000000",
        20 => "11111101111010000000000000001100",
        21 => "11111001000000000000110000000000",
        22 => "11110000000000000000000000000001",
        23 => "11111101110000000000101010000000",
        24 => "11111101111010000000000000001100",
        25 => "11111001000000000000110000000000",
        26 => "11110000100000000000000000000001",
        27 => "11110110011000000000000000001001",
        others => (others => '0')
    );