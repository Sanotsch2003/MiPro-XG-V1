    signal ram : ram_type :=(
        0 => "11110110110000000000000000000110",
        1 => "11111101110000000001011111000000",
        2 => "11111101110000000001011111000001",
        3 => "11111101110000000010101010000010",
        4 => "11111101110000000001111000000011",
        5 => "11110110110000000000000000001100",
        6 => "11110100001000000000000000000000",
        7 => "11111101110000000000000000001001",
        8 => "11111101111100000000000000001100",
        9 => "11111001000000000000110010011001",
        10 => "11111101110000000000000000001010",
        11 => "11111101110100101100000000001011",
        12 => "11111011100000000000101110011011",
        13 => "11110000100000000000000010011010",
        14 => "11111011110000000000100101001001",
        15 => "11111010101000000000100110110000",
        16 => "00010110011000000000000000000100",
        17 => "11111101100000000000000110101111",
        18 => "11111101110000000000000000001010",
        19 => "11111101111100000000000000001100",
        20 => "11111001000000000000110010101010",
        21 => "11111101110000000000101000001100",
        22 => "11111110000000000000000011001011",
        23 => "11111011100000000000101010111000",
        24 => "11111110000000000000000111001011",
        25 => "11111011100000000000101010111010",
        26 => "11111101110000000000100110001100",
        27 => "11111011100000000000101011001010",
        28 => "11111101110000000000110010001011",
        29 => "11111101110000000000101000001100",
        30 => "11111110000000000000101111001011",
        31 => "11111011100000000000101110101011",
        32 => "11111101110111111111111111101001",
        33 => "11111101100010100000000100100111",
        34 => "11110000100000000000000010001001",
        35 => "11110000100000000000000010100111",
        36 => "11111011100000000000101011001010",
        37 => "11111011100000000000100011001000",
        38 => "11111010101000000000101010110000",
        39 => "00010110011000000000000000000110",
        40 => "11111101100000000000000110101111",
        others => (others => '0')
    );