    signal ram : ram_type :=(
        0 => "11111101110000000000101000000000",
        1 => "11111101111010000000000000001100",
        2 => "11111001000000000000110000000000",
        3 => "11111101110001001000010010000001",
        4 => "11111101111000000001111010001100",
        5 => "11111001000000000000110000010001",
        6 => "11110000100000000000000000000001",
        7 => "11111101110000000000101010000000",
        8 => "11111101111010000000000000001100",
        9 => "11111001000000000000110000000000",
        10 => "11111101110000000000000010100001",
        11 => "11111101110000000000000000000010",
        12 => "11110000100000000000000000000010",
        13 => "11111101110000000000000000000011",
        14 => "11111011110000000000001100010011",
        15 => "11111010101000000000001100010000",
        16 => "00010110011000000000000000000011",
        17 => "11111011110000000000001000010010",
        18 => "11110110011000000000000000000111",
        others => (others => '0')
    );