    signal ram : ram_type :=(
        0 => "11111101110010101010101010100000",
        1 => "11111101111010101010101010101100",
        2 => "11111001000000000000110000000000",
        others => (others => '0')
    );