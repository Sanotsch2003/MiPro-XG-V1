    signal ram : ram_type :=(
        0 => "11111101110111111100000000000000",
        1 => "11111101111001111111111111101100",
        2 => "11111001000000000000110000000000",
        3 => "11111101110000000001111010000001",
        4 => "11111101111000000000000000001100",
        5 => "11111001000000000000110000010001",
        6 => "11110000100000000000000000000001",
        7 => "11111101110111111100000010000000",
        8 => "11111101111001111111111111101100",
        9 => "11111001000000000000110000000000",
        10 => "11111101110000000000000000100001",
        11 => "11110000100000000000000000000001",
        12 => "11111101110111111100000100000000",
        13 => "11111101111001111111111111101100",
        14 => "11111001000000000000110000000000",
        15 => "11111101110000000010010100000001",
        16 => "11111101111000000000000000001100",
        17 => "11111001000000000000110000010001",
        18 => "11110000100000000000000000000001",
        19 => "11111101110111111100000110000000",
        20 => "11111101111001111111111111101100",
        21 => "11111001000000000000110000000000",
        22 => "11111101110000000000000000100001",
        23 => "11110000100000000000000000000001",
        24 => "11111101110111111100001000000000",
        25 => "11111101111001111111111111101100",
        26 => "11111001000000000000110000000000",
        27 => "11111101110000000010101110000001",
        28 => "11111101111000000000000000001100",
        29 => "11111001000000000000110000010001",
        30 => "11110000100000000000000000000001",
        31 => "11111101110111111100001010000000",
        32 => "11111101111001111111111111101100",
        33 => "11111001000000000000110000000000",
        34 => "11111101110000000000000000100001",
        35 => "11110000100000000000000000000001",
        36 => "11111101110111111100001100000000",
        37 => "11111101111001111111111111101100",
        38 => "11111001000000000000110000000000",
        39 => "11111101110000000011001000000001",
        40 => "11111101111000000000000000001100",
        41 => "11111001000000000000110000010001",
        42 => "11110000100000000000000000000001",
        43 => "11111101110111111100001110000000",
        44 => "11111101111001111111111111101100",
        45 => "11111001000000000000110000000000",
        46 => "11111101110000000000000000100001",
        47 => "11110000100000000000000000000001",
        48 => "11111101110111111100011100000000",
        49 => "11111101111001111111111111101100",
        50 => "11111001000000000000110000000000",
        51 => "11111101110000000011100010000001",
        52 => "11111101111000000000000000001100",
        53 => "11111001000000000000110000010001",
        54 => "11110000100000000000000000000001",
        55 => "11111101110111111100011110000000",
        56 => "11111101111001111111111111101100",
        57 => "11111001000000000000110000000000",
        58 => "11111101110000000000000000100001",
        59 => "11110000100000000000000000000001",
        60 => "11110110010000000000000000111010",
        61 => "11111101110000000000101000000000",
        62 => "11111101111010000000000000001100",
        63 => "11111001000000000000110000000000",
        64 => "11111101110001001000011010000001",
        65 => "11111101111000000001111010001100",
        66 => "11111001000000000000110000010001",
        67 => "11110000100000000000000000000001",
        68 => "11111101110000000000101010000000",
        69 => "11111101111010000000000000001100",
        70 => "11111001000000000000110000000000",
        71 => "11111101110111011100000000000001",
        72 => "11110000100000000000000000000001",
        73 => "11110100001000000000000000000000",
        74 => "11111101110000000000101000000000",
        75 => "11111101111010000000000000001100",
        76 => "11111001000000000000110000000000",
        77 => "11111101110001001000011010000001",
        78 => "11111101111000000001111010001100",
        79 => "11111001000000000000110000010001",
        80 => "11110000100000000000000000000001",
        81 => "11111101110000000000101010000000",
        82 => "11111101111010000000000000001100",
        83 => "11111001000000000000110000000000",
        84 => "11111101110111011100000000100001",
        85 => "11110000100000000000000000000001",
        86 => "11110100001000000000000000000000",
        87 => "11111101110000000000101000000000",
        88 => "11111101111010000000000000001100",
        89 => "11111001000000000000110000000000",
        90 => "11111101110001001000011010000001",
        91 => "11111101111000000001111010001100",
        92 => "11111001000000000000110000010001",
        93 => "11110000100000000000000000000001",
        94 => "11111101110000000000101010000000",
        95 => "11111101111010000000000000001100",
        96 => "11111001000000000000110000000000",
        97 => "11111101110111011100000001000001",
        98 => "11110000100000000000000000000001",
        99 => "11110100001000000000000000000000",
        100 => "11111101110000000000101000000000",
        101 => "11111101111010000000000000001100",
        102 => "11111001000000000000110000000000",
        103 => "11111101110001001000011010000001",
        104 => "11111101111000000001111010001100",
        105 => "11111001000000000000110000010001",
        106 => "11110000100000000000000000000001",
        107 => "11111101110000000000101010000000",
        108 => "11111101111010000000000000001100",
        109 => "11111001000000000000110000000000",
        110 => "11111101110111011100000001100001",
        111 => "11110000100000000000000000000001",
        112 => "11110100001000000000000000000000",
        113 => "11111011110000000000011000010110",
        114 => "11111101110000000000101010000111",
        115 => "11111101111010000000000000001100",
        116 => "11111001000000000000110001110111",
        117 => "11110000100000000000000001110110",
        118 => "11110100100000000000000000000000",
        119 => "11111101110000000000101000000000",
        120 => "11111101111010000000000000001100",
        121 => "11111001000000000000110000000000",
        122 => "11111101110001001000010010000001",
        123 => "11111101111000000001111010001100",
        124 => "11111001000000000000110000010001",
        125 => "11110000100000000000000000000001",
        126 => "11111101110000000001001110000000",
        127 => "11111101111010000000000000001100",
        128 => "11111001000000000000110000000000",
        129 => "11111101110111100001000000000001",
        130 => "11111101111000000101111101001100",
        131 => "11111001000000000000110000010001",
        132 => "11110000100000000000000000000001",
        133 => "11111101110000000001010000000000",
        134 => "11111101111010000000000000001100",
        135 => "11111001000000000000110000000000",
        136 => "11111101110000000000000001100001",
        137 => "11110000100000000000000000000001",
        138 => "11111101110000000000111000000000",
        139 => "11111101111010000000000000001100",
        140 => "11111001000000000000110000000000",
        141 => "11111101110000000000000000100001",
        142 => "11110000100000000000000000000001",
        143 => "11111101110000000001010100000000",
        144 => "11111101111010000000000000001100",
        145 => "11111001000000000000110000000000",
        146 => "11111101110000000000000001000001",
        147 => "11110000100000000000000000000001",
        148 => "11111101110000000001011100000000",
        149 => "11111101111010000000000000001100",
        150 => "11111001000000000000110000000000",
        151 => "11111101110000000000000001000001",
        152 => "11110000100000000000000000000001",
        153 => "11111101110000000001100100000000",
        154 => "11111101111010000000000000001100",
        155 => "11111001000000000000110000000000",
        156 => "11111101110000000000000001000001",
        157 => "11110000100000000000000000000001",
        158 => "11111101110000000001011000000000",
        159 => "11111101111010000000000000001100",
        160 => "11111001000000000000110000000000",
        161 => "11111101110000000001100000000001",
        162 => "11111101111010000000000000001100",
        163 => "11111001000000000000110000010001",
        164 => "11111101110000000001101000000010",
        165 => "11111101111010000000000000001100",
        166 => "11111001000000000000110000100010",
        167 => "11111101110000000001111111100011",
        168 => "11111101110000000000000000000100",
        169 => "11111101110000000000000000000101",
        170 => "11110110110000000000000000011001",
        171 => "11110110110000000000000000010010",
        172 => "11110110110000000000000000010111",
        173 => "11111010110000000000001100010011",
        174 => "11111011110000000000010000010100",
        175 => "11111010111000000000001100000000",
        176 => "00010110011000000000000000000110",
        177 => "11110110110000000000000000001100",
        178 => "11110110110000000000000000010001",
        179 => "11111010110000000000010000010100",
        180 => "11111011110000000000010100010101",
        181 => "11111010111000000000010000000000",
        182 => "00010110011000000000000000000110",
        183 => "11110110110000000000000000000110",
        184 => "11110110110000000000000000001011",
        185 => "11111010110000000000010100010101",
        186 => "11111011110000000000001100010011",
        187 => "11111010111000000000010100000000",
        188 => "00010110011000000000000000000110",
        189 => "11110110011000000000000000010011",
        190 => "11111101110000000000000000001010",
        191 => "11111101110011101010011000001011",
        192 => "11111010101000000000101110100000",
        193 => "00001101100000000000000110101111",
        194 => "11111011110000000000101000011010",
        195 => "11110110011000000000000000000100",
        196 => "11110000100000000000000000000011",
        197 => "11110000100000000000000000010100",
        198 => "11110000100000000000000000100101",
        199 => "11111101100000000000000110101111",
        others => (others => '0')
    );