library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity CPU_Core is
    Generic(
        numInterrupts : integer := 5
    );

    Port (
        enable                  : in std_logic;
        hardwareReset           : in std_logic;
        clk                     : in std_logic;
        alteredClock            : in std_logic;

        programmingMode         : in std_logic;

        dataIn                  : in std_logic_vector(31 downto 0);
        dataOut                 : out std_logic_vector(31 downto 0);
        addressOut              : out std_logic_vector(31 downto 0);
        
        readEn                  : out std_logic;
        writeEn                 : out std_logic;
        softwareReset           : out std_logic;
        memOpFinished           : in std_logic;

        --interupt vector table and interrupt priority register
        IVT                     : in std_logic_vector(numInterrupts*32-1 downto 0);
        PR                      : in std_logic_vector(numInterrupts*3-1 downto 0);

        externalInterrupts      : in std_logic_vector(numInterrupts-1 downto 0); --there are no internal interrupts so far
        clearExternalInterrupts : out std_logic_vector(numInterrupts-1 downto 0); 

        --debugging
        debug                   : out std_logic_vector(866+numInterrupts-1 downto 0)
    );
end CPU_Core;

architecture Behavioral of CPU_Core is
    component ALU is
        port (
            operand1             : in std_logic_vector(31 downto 0);
            operand2             : in std_logic_vector(31 downto 0);
    
            bitManipulationCode  : in std_logic_vector(1 downto 0);
            bitManipulationValue : in std_logic_vector(4 downto 0);
    
            opCode               : in std_logic_vector(3 downto 0);
            carryIn              : in std_logic;
            
            upperSel             : in std_logic;
    
            --outputs
            result               : out std_logic_vector(31 downto 0);
            flagsCPSR            : out std_logic_vector(3 downto 0);
            debug                : out std_logic_vector(99 downto 0)   
         );
    end component;

    component registerFile is
        port(
            enable           : in std_logic;
            reset            : in std_logic;
            clk              : in std_logic;
            alteredClock     : in std_logic;
    
            dataIn           : in std_logic_vector(31 downto 0);
            loadRegistersSel : in std_logic_vector(15 downto 0);
            dataOut          : out std_logic_vector(16 * 32-1 downto 0)
        );
    end component;

    component busManagement is
        Port ( 
              dataFromRegisters   : in std_logic_vector(16 * 32-1 downto 0);
              dataFromCU          : in std_logic_vector(31 downto 0);
              dataFromALU         : in std_logic_vector(31 downto 0);
              dataFromMem         : in std_logic_vector(31 downto 0);
      
              operand1            : out std_logic_vector(31 downto 0);
              operand2            : out std_logic_vector(31 downto 0);
      
              operand1Sel         : in std_logic_vector(4 downto 0);
              operand2Sel         : in std_logic_vector(4 downto 0); 
      
              dataToRegisters     : out std_logic_vector(31 downto 0);
      
              dataToRegistersSel  : in std_logic
        );
    end component;

    component coreInterruptController is
        Generic(
            numInterrupts : integer := 5
          );
          Port (
            interruptSignals : in std_logic_vector(numInterrupts-1 downto 0);
        
            IVT_in           : in std_logic_vector(32 * numInterrupts - 1 downto 0);
            PR_in            : in std_logic_vector(3 * numInterrupts - 1 downto 0);
        
            vectorOut        : out std_logic_vector(31 downto 0)
           );
    end component;

    component controlUnit is
        Generic(
            numInterrupts : integer := 5
        );
        Port(
            enable              : in std_logic;
            hardwareReset       : in std_logic;
            softwareReset       : out std_logic;
            clk                 : in std_logic;
            alteredClock        : in std_logic;
    
            --control signals generated by CU
            operand1Sel         : out std_logic_vector(4 downto 0);
            operand2Sel         : out std_logic_vector(4 downto 0); 
    
            dataToRegistersSel  : out std_logic;
            loadRegistersSel    : out std_logic_vector(15 downto 0);
    
            bitManipulationCode : out std_logic_vector(1 downto 0);
            bitManipulationValue: out std_logic_vector(4 downto 0);
    
            opCode              : out std_logic_vector(3 downto 0);
            carryIn             : out std_logic;
            upperSel            : out std_logic;
    
            clearInterrupts     : out std_logic_vector(numInterrupts-1 downto 0);
              
            --signals controlling the CU
            programmingMode     : in std_logic;
            IVT_address         : in std_logic_vector(31 downto 0);
            PC                  : in std_logic_vector(31 downto 0);
            flagsCPSR           : in std_logic_vector(3 downto 0);
            memOpFinished       : in std_logic;
    
            --debug signals
            debug : out std_logic_vector(49 downto 0)
    );
    end component;

    --internal signals
    --ALU
    signal operand1 : std_logic_vector(31 downto 0);
    signal operand2 : std_logic_vector(31 downto 0);
    signal bitManipulationCode : std_logic_vector(1 downto 0);
    signal bitManipulationValue : std_logic_vector(4 downto 0);
    signal opCode : std_logic_vector(3 downto 0);
    signal carryIn : std_logic;
    signal upperSel : std_logic;
    
    --register file
    signal dataToRegisters  : std_logic_vector(31 downto 0);
    signal loadRegistersSel : std_logic_vector(15 downto 0);

    --bus management
    signal dataFromRegisters   : std_logic_vector(16 * 32-1 downto 0);
    signal dataFromCU          : std_logic_vector(31 downto 0);
    signal dataFromALU         : std_logic_vector(31 downto 0);
    signal dataFromMem         : std_logic_vector(31 downto 0);
    signal operand1Sel         : std_logic_vector(4 downto 0);
    signal operand2Sel         : std_logic_vector(4 downto 0); 
    signal dataToRegistersSel  : std_logic;

    --interrupt controller
    --signal internalInterrupts  --should be uncommented if any internal interrupts are being used
    signal interrupts               : std_logic_vector(numInterrupts-1 downto 0);
    signal interruptHandlerAddress  : std_logic_vector(31 downto 0);
    --signal clearInternalInterrupts --should be uncommented if any internal interrupts are being used
    signal clearInterrupts          : std_logic_vector(numInterrupts-1 downto 0);

    --CU
    signal ALU_flags  : std_logic_vector(3 downto 0);

    --debug signals
    signal ALU_debug : std_logic_vector(99 downto 0);
    signal CU_debug  : std_logic_vector(49 downto 0);

    --others
    signal reset               : std_logic;
    signal softwareResetFromCu : std_logic;

begin
    --reset signals
    reset <= hardwareReset or softwareResetFromCu;
    softwareReset <= softwareResetFromCu;

    --data signals
    dataFromMem <= dataIn;

    --interrupts
    --interrupts <= internalInterrupts & externalInterrupts -- if any internal interrupts are being used
    interrupts              <= externalInterrupts;
    clearExternalInterrupts <= clearInterrupts; --when internal interrupts are used only the external once should be passed to the clearExternalInterrupts signal

    --       32 bit        4 bit       100 bit     512 bit             32 bit     32 bit     32 bit            32 Bit                    5 Bit         5 Bit         1 Bit                16 Bit             2 Bit                 5 Bit                  3 Bit    1 Bit     1 Bit      1 Bit                 numInterrupts Bit 50 Bit
    debug <= dataFromALU & ALU_flags & ALU_debug & dataFromRegisters & operand1 & operand2 & dataToRegisters & interruptHandlerAddress & operand1Sel & operand2Sel & dataToRegistersSel & loadRegistersSel & bitManipulationCode & bitManipulationValue & opCode & carryIn & upperSel & softwareResetFromCu & clearInterrupts & CU_debug;

    ALU_inst : ALU
        port map(
            --inputs
            operand1                => operand1,          
            operand2                => operand2,             
    
            bitManipulationCode     => bitManipulationCode,
            bitManipulationValue    => bitManipulationValue,
    
            opCode                  => opCode,
            carryIn                 => carryIn,
            
            upperSel                => upperSel,        
    
            --outputs
            result                  => dataFromALU,
            flagsCPSR               => ALU_flags,
            debug                   => ALU_debug
        );

    RegisterFile_inst : registerFile
        port map(
            --inputs
            enable              => enable,     
            reset               => reset,
            clk                 => clk,
            alteredClock        => alteredClock,
    
            dataIn              => dataToRegisters,
            loadRegistersSel    => loadRegistersSel,
            --output
            dataOut             => dataFromRegisters
        );

    busManagement_inst : busManagement
        port map(
            --inputs
            dataFromRegisters       => dataFromRegisters,
            dataFromCU              => dataFromCU,
            dataFromALU             => dataFromALU,
            dataFromMem             => dataFromMeM,
      
            operand1Sel             => operand1Sel,
            operand2Sel             => operand2Sel,

            dataToRegistersSel      => dataToRegistersSel,

            --outputs
            operand1                => operand1,            
            operand2                => operand2,
            dataToRegisters         => dataToRegisters
      
        );

    interruptControler_inst : coreInterruptController
        generic map(
            numInterrupts => numInterrupts
        )
        port map(
            --inputs
            interruptSignals => interrupts,
            IVT_in           => IVT, 
            PR_in            => PR,
            --output
            vectorOut        => interruptHandlerAddress
        );

    CU : controlUnit
        generic map(
            numInterrupts => numInterrupts
        )
        port map(
            --inputs
            enable                  => enable,
            hardwareReset           => hardwareReset,
            clk                     => clk,
            alteredClock            => alteredClock,

            programmingMode         => programmingMode,
            IVT_address             => interruptHandlerAddress,
            PC                      => dataFromRegisters(16*32-1 downto 15*32), --program counter
            flagsCPSR               => ALU_flags,
            memOpFinished           => memOpFinished,

            --outputs
            operand1Sel             => operand1Sel,
            operand2Sel             => operand2Sel,
    
            dataToRegistersSel      => dataToRegistersSel,
            loadRegistersSel        => loadRegistersSel,
    
            bitManipulationCode     => bitManipulationCode,
            bitManipulationValue    => bitManipulationValue,
    
            opCode                  => opCode,
            carryIn                 => carryIn,
            upperSel                => upperSel,

            softwareReset           => softwareResetFromCu,
            clearInterrupts         => clearInterrupts,
              
            debug                   => CU_debug
        );
        

end Behavioral;
