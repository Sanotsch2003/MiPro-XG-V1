    signal ram : ram_type :=(
        0 => "11111101110000000000101000000000",
        1 => "11111101111010000000000000001100",
        2 => "11111001000000000000110000000000",
        3 => "11111101110001001000010001100001",
        4 => "11111101111000000001111010001100",
        5 => "11111001000000000000110000010001",
        6 => "11110000100000000000000000000001",
        7 => "11111011110000000000111101001101",
        8 => "11110110110000000000000000000100",
        9 => "11111011110000000000011100010111",
        10 => "11111011110000000000111101001101",
        11 => "11110110110000000000000000000110",
        12 => "11110110011000000000000000000110",
        13 => "11111101110000000000101010001011",
        14 => "11111101111010000000000000001100",
        15 => "11111001000000000000110010111011",
        16 => "11110000100000000000000010110111",
        17 => "11111101100000000000000110101111",
        18 => "11111101110000000000000000001010",
        19 => "11111101110111000110110000001011",
        20 => "11111101111000000000001011001100",
        21 => "11111001000000000000110010111011",
        22 => "11111010101000000000101110100000",
        23 => "00001101100000000000000110101111",
        24 => "11111011110000000000101000011010",
        25 => "11110110011000000000000000000100",
        others => (others => '0')
    );