LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY CPU_Core IS
    GENERIC (
        numExternalInterrupts   : INTEGER;
        numInterrupts           : INTEGER;
        numCPU_CoreDebugSignals : INTEGER
    );
    PORT (
        enable     : IN STD_LOGIC;
        reset      : IN STD_LOGIC;
        clk        : IN STD_LOGIC;
        alteredClk : IN STD_LOGIC;

        programmingMode : IN STD_LOGIC;

        dataFromMem : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        dataOut     : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
        addressOut  : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);

        memWriteReq   : OUT STD_LOGIC;
        memReadReq    : OUT STD_LOGIC;
        softwareReset : OUT STD_LOGIC;
        memOpFinished : IN STD_LOGIC;

        --interupt vector table and interrupt priority register
        IVT : IN STD_LOGIC_VECTOR(numInterrupts * 32 - 1 DOWNTO 0);
        IPR : IN STD_LOGIC_VECTOR(numInterrupts * 3 - 1 DOWNTO 0);

        externalInterrupts    : IN STD_LOGIC_VECTOR(numExternalInterrupts - 1 DOWNTO 0); --there are no internal interrupts so far
        externalInterruptsClr : OUT STD_LOGIC_VECTOR(numExternalInterrupts - 1 DOWNTO 0);

        --debugging
        debug : OUT STD_LOGIC_VECTOR(numCPU_CoreDebugSignals - 1 DOWNTO 0)
    );
END CPU_Core;

ARCHITECTURE Behavioral OF CPU_Core IS
    COMPONENT ALU IS
        PORT (
            clk        : IN STD_LOGIC;
            reset      : IN STD_LOGIC;
            enable     : IN STD_LOGIC;
            alteredClk : IN STD_LOGIC;
            operand1   : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
            operand2   : IN STD_LOGIC_VECTOR(31 DOWNTO 0);

            bitManipulationCode  : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
            bitManipulationValue : IN STD_LOGIC_VECTOR(4 DOWNTO 0);

            opCode  : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
            carryIn : IN STD_LOGIC;

            upperSel : IN STD_LOGIC;

            --outputs
            result    : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
            flagsCPSR : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
            debug     : OUT STD_LOGIC_VECTOR(67 DOWNTO 0)
        );
    END COMPONENT;

    COMPONENT registerFile IS
        PORT (
            enable     : IN STD_LOGIC;
            reset      : IN STD_LOGIC;
            clk        : IN STD_LOGIC;
            alteredClk : IN STD_LOGIC;

            dataIn           : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
            loadRegistersSel : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
            dataOut          : OUT STD_LOGIC_VECTOR(16 * 32 - 1 DOWNTO 0);
            createLink       : IN STD_LOGIC
        );
    END COMPONENT;

    COMPONENT busManagement IS
        PORT (
            dataFromRegisters          : IN STD_LOGIC_VECTOR(16 * 32 - 1 DOWNTO 0);
            dataFromCU                 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
            dataFromALU                : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
            dataFromMem                : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
            bitManipulationValueFromCU : IN STD_LOGIC_VECTOR(4 DOWNTO 0);

            operand1              : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
            operand2              : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
            dataToMem             : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
            bitManipulationValOut : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);

            operand1Sel           : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
            operand2Sel           : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
            dataToMemSel          : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
            bitManipulationValSel : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
            dataToRegisters       : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
            dataToRegistersSel    : IN STD_LOGIC
        );
    END COMPONENT;

    COMPONENT coreInterruptController IS
        GENERIC (
            numInterrupts : INTEGER
        );
        PORT (
            clk        : IN STD_LOGIC;
            interrupts : IN STD_LOGIC_VECTOR(numInterrupts - 1 DOWNTO 0);

            IVT_in : IN STD_LOGIC_VECTOR(32 * numInterrupts - 1 DOWNTO 0);
            IPR_in : IN STD_LOGIC_VECTOR(3 * numInterrupts - 1 DOWNTO 0);

            interruptIndex          : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            interruptHandlerAddress : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
        );
    END COMPONENT;

    COMPONENT controlUnit IS
        GENERIC (
            numInterrupts : INTEGER := 10
        );

        PORT (
            enable        : IN STD_LOGIC;
            reset         : IN STD_LOGIC;
            softwareReset : OUT STD_LOGIC;
            clk           : IN STD_LOGIC;
            alteredClk    : IN STD_LOGIC;

            --control signals generated by CU
            operand1Sel  : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
            operand2Sel  : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
            dataToMemSel : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);

            dataToRegistersSel    : OUT STD_LOGIC;
            loadRegistersSel      : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
            createLink            : OUT STD_LOGIC;
            bitManipulationValSel : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);

            bitManipulationCode  : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
            bitManipulationValue : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);

            ALU_opCode : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
            carryIn    : OUT STD_LOGIC;
            upperSel   : OUT STD_LOGIC;

            memWriteReq : OUT STD_LOGIC;
            memReadReq  : OUT STD_LOGIC;

            interruptsClr : OUT STD_LOGIC_VECTOR(numInterrupts - 3 DOWNTO 0);
            dataToALU     : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);

            ALU_En : OUT STD_LOGIC;

            --Interrupt signals
            interrupts : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);

            --signals controlling the CU
            PC                      : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
            programmingMode         : IN STD_LOGIC;
            InterruptHandlerAddress : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
            interruptIndex          : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
            dataFromMem             : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
            dataFromALU             : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
            flagsFromALU            : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
            memOpFinished           : IN STD_LOGIC;
            --debug signals
            debug : OUT STD_LOGIC_VECTOR(38 DOWNTO 0)
        );
    END COMPONENT;

    --internal signals
    --ALU
    SIGNAL ALU_En               : STD_LOGIC;
    SIGNAL operand1             : STD_LOGIC_VECTOR(31 DOWNTO 0);
    SIGNAL operand2             : STD_LOGIC_VECTOR(31 DOWNTO 0);
    SIGNAL bitManipulationCode  : STD_LOGIC_VECTOR(1 DOWNTO 0);
    SIGNAL bitManipulationValue : STD_LOGIC_VECTOR(4 DOWNTO 0);
    SIGNAL ALU_opCode           : STD_LOGIC_VECTOR(3 DOWNTO 0);
    SIGNAL carryIn              : STD_LOGIC;
    SIGNAL upperSel             : STD_LOGIC;

    --register file
    SIGNAL dataToRegisters  : STD_LOGIC_VECTOR(31 DOWNTO 0);
    SIGNAL loadRegistersSel : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL createLink       : STD_LOGIC;

    --bus management
    SIGNAL dataFromRegisters          : STD_LOGIC_VECTOR(16 * 32 - 1 DOWNTO 0);
    SIGNAL dataFromCU                 : STD_LOGIC_VECTOR(31 DOWNTO 0);
    SIGNAL dataFromALU                : STD_LOGIC_VECTOR(31 DOWNTO 0);
    SIGNAL operand1Sel                : STD_LOGIC_VECTOR(4 DOWNTO 0);
    SIGNAL operand2Sel                : STD_LOGIC_VECTOR(4 DOWNTO 0);
    SIGNAL dataToMemSel               : STD_LOGIC_VECTOR(3 DOWNTO 0);
    SIGNAL dataToRegistersSel         : STD_LOGIC;
    SIGNAL bitManipulationValSel      : STD_LOGIC_VECTOR(4 DOWNTO 0);
    SIGNAL bitManipulationValueFromCU : STD_LOGIC_VECTOR(4 DOWNTO 0);

    --interrupt controller
    --signal internalInterrupts  --should be uncommented if any internal interrupts are being used
    SIGNAL interrupts              : STD_LOGIC_VECTOR(numInterrupts - 1 DOWNTO 0);
    SIGNAL interruptHandlerAddress : STD_LOGIC_VECTOR(31 DOWNTO 0);
    SIGNAL interruptIndex          : STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL interruptsClr           : STD_LOGIC_VECTOR(numInterrupts - 3 DOWNTO 0);

    --CU
    SIGNAL ALU_flags     : STD_LOGIC_VECTOR(3 DOWNTO 0);
    SIGNAL ALU_EnFromCU  : STD_LOGIC;
    SIGNAL CU_interrupts : STD_LOGIC_VECTOR(1 DOWNTO 0);

    --debug signals
    SIGNAL ALU_debug : STD_LOGIC_VECTOR(67 DOWNTO 0);
    SIGNAL CU_debug  : STD_LOGIC_VECTOR(38 DOWNTO 0);

    --output signals
    SIGNAL dataToMem      : STD_LOGIC_VECTOR(31 DOWNTO 0);
    SIGNAL CU_memWriteReq : STD_LOGIC;
    SIGNAL CU_memReadReq  : STD_LOGIC;

BEGIN
    --enable signals
    ALU_En <= enable AND ALU_EnFromCU;

    --interrupts
    interrupts            <= externalInterrupts & CU_interrupts;
    externalInterruptsClr <= interruptsClr(numInterrupts - 3 DOWNTO numInterrupts - 2 - numExternalInterrupts);

    --assigning output signals
    memWriteReq <= CU_memWriteReq;
    memReadReq  <= CU_memReadReq;
    dataOut     <= dataToMem;
    addressOut  <= dataFromALU;

    ---             32 Bit        4 Bit       68 Bit      32 Bit       512 Bit             32 Bit     32 Bit     32 Bit      32 Bit        5 Bit         5 Bit         1 Bit                16 Bit             2 Bit                 5 Bit                  3 Bit        1 Bit     1 Bit      1 Bit numInterrupts Bit 38 Bit     1Bit             1 Bit        
    debug <= dataFromALU & ALU_flags & ALU_debug & dataFromCU & dataFromRegisters & operand1 & operand2 & dataToMem & dataFromMem & operand1Sel & operand2Sel & dataToRegistersSel & loadRegistersSel & bitManipulationCode & bitManipulationValue & ALU_opCode & carryIn & upperSel & '0' & "0000000000" & CU_debug & CU_memWriteReq & CU_memReadReq;
    --debug <= (others => '0');

    ALU_inst : ALU
    PORT MAP(
        --inputs
        clk        => clk,
        reset      => reset,
        enable     => ALU_En,
        alteredClk => alteredClk,
        operand1   => operand1,
        operand2   => operand2,

        bitManipulationCode  => bitManipulationCode,
        bitManipulationValue => bitManipulationValue,

        opCode  => ALU_opCode,
        carryIn => carryIn,

        upperSel => upperSel,

        --outputs
        result    => dataFromALU,
        flagsCPSR => ALU_flags,
        debug     => ALU_debug
    );

    RegisterFile_inst : registerFile
    PORT MAP(
        --inputs
        enable     => enable,
        reset      => reset,
        clk        => clk,
        alteredClk => alteredClk,

        dataIn           => dataToRegisters,
        loadRegistersSel => loadRegistersSel,
        createLink       => createLink,
        --output
        dataOut => dataFromRegisters
    );

    busManagement_inst : busManagement
    PORT MAP(
        --inputs    
        dataFromRegisters          => dataFromRegisters,
        dataFromCU                 => dataFromCU,
        dataFromALU                => dataFromALU,
        dataFromMem                => dataFromMeM,
        bitManipulationValueFromCU => bitManipulationValueFromCU,

        operand1Sel           => operand1Sel,
        operand2Sel           => operand2Sel,
        dataToMemSel          => dataToMemSel,
        bitManipulationValSel => bitManipulationValSel,

        dataToRegistersSel => dataToRegistersSel,

        --outputs
        operand1              => operand1,
        operand2              => operand2,
        dataToMem             => dataToMem,
        dataToRegisters       => dataToRegisters,
        bitManipulationValOut => bitManipulationValue
    );

    interruptController_inst : coreInterruptController
    GENERIC MAP(
        numInterrupts => numInterrupts
    )
    PORT MAP(
        --inputs
        clk        => clk,
        interrupts => interrupts,
        IVT_in     => IVT,
        IPR_in     => IPR,
        --output
        interruptHandlerAddress => interruptHandlerAddress,
        interruptIndex          => interruptIndex
    );

    CU : controlUnit
    GENERIC MAP(
        numInterrupts => numInterrupts
    )
    PORT MAP(
        --inputs
        enable     => enable,
        reset      => reset,
        clk        => clk,
        alteredClk => alteredClk,

        programmingMode         => programmingMode,
        interruptHandlerAddress => interruptHandlerAddress,
        interruptIndex          => interruptIndex,
        dataFromMem             => dataFromMem,
        dataFromALU             => dataFromALU,
        flagsFromALU            => ALU_flags,
        memOpFinished           => memOpFinished,
        PC                      => dataFromRegisters(16 * 32 - 1 DOWNTO 15 * 32),

        --outputs
        operand1Sel  => operand1Sel,
        operand2Sel  => operand2Sel,
        dataToMemSel => dataToMemSel,

        dataToRegistersSel    => dataToRegistersSel,
        createLink            => createLink,
        loadRegistersSel      => loadRegistersSel,
        bitManipulationValSel => bitManipulationValSel,

        bitManipulationCode  => bitManipulationCode,
        bitManipulationValue => bitManipulationValueFromCU,

        ALU_opCode => ALU_opCode,
        ALU_En     => ALU_EnFromCU,
        carryIn    => carryIn,
        upperSel   => upperSel,

        memWriteReq => CU_memWriteReq,
        memReadReq  => CU_memReadReq,

        softwareReset => softwareReset,
        interruptsClr => interruptsClr,

        dataToALU => dataFromCU,

        interrupts => CU_interrupts,

        debug => CU_debug
    );
END Behavioral;