    signal ram : ram_type :=(
        0 => "11110000",
        1 => "00111010",
        2 => "10101011",
        3 => "11101111",
        others => (others => '0')
    );