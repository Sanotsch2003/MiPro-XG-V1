    signal ram : ram_type :=(
        0 => "11111101110000000000101000000000",
        1 => "11111101111010000000000000001100",
        2 => "11111001000000000000110000000000",
        3 => "11111101110001001000010010000001",
        4 => "11111101111000000001111010001100",
        5 => "11111001000000000000110000010001",
        6 => "11110000100000000000000000000001",
        7 => "11110110110000000000000000000011",
        8 => "11111011110000000000011100010111",
        9 => "11110110110000000000000000000110",
        10 => "11110110011000000000000000000100",
        11 => "11111101110000000000101010001011",
        12 => "11111101111010000000000000001100",
        13 => "11111001000000000000110010111011",
        14 => "11110000100000000000000010110111",
        15 => "11111101100000000000000110101111",
        16 => "11111101110000000000000000001010",
        17 => "11111101110111000110110000001011",
        18 => "11111101111000000000001011001100",
        19 => "11111001000000000000110010111011",
        20 => "11111010101000000000101110100000",
        21 => "00001101100000000000000110101111",
        22 => "11111011110000000000101000011010",
        23 => "11110110011000000000000000000100",
        others => (others => '0')
    );