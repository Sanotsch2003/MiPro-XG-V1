LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

--TODO operandXSel <= operandXSelReg is conditionally assigned. should also work if it is always assigned

ENTITY controlUnit IS
    GENERIC (
        numInterrupts : INTEGER := 10
    );

    PORT (
        enable        : IN STD_LOGIC;
        reset         : IN STD_LOGIC;
        softwareReset : OUT STD_LOGIC;
        clk           : IN STD_LOGIC;
        alteredClk    : IN STD_LOGIC;

        --control signals generated by CU
        operand1Sel  : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
        operand2Sel  : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
        dataToMemSel : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);

        dataToRegistersSel    : OUT STD_LOGIC;
        loadRegistersSel      : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
        createLink            : OUT STD_LOGIC;
        bitManipulationValSel : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);

        bitManipulationCode  : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
        bitManipulationValue : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);

        ALU_opCode : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
        carryIn    : OUT STD_LOGIC;
        upperSel   : OUT STD_LOGIC;

        memWriteReq : OUT STD_LOGIC;
        memReadReq  : OUT STD_LOGIC;

        interruptsClr : OUT STD_LOGIC_VECTOR(numInterrupts - 3 DOWNTO 0);
        dataToALU     : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);

        ALU_En : OUT STD_LOGIC;

        --Interrupt signals
        interrupts : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);

        --signals controlling the CU
        PC                      : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        programmingMode         : IN STD_LOGIC;
        InterruptHandlerAddress : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        interruptIndex          : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
        dataFromMem             : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        dataFromALU             : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        flagsFromALU            : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        memOpFinished           : IN STD_LOGIC;
        --debug signals
        debug : OUT STD_LOGIC_VECTOR(38 DOWNTO 0)
    );
END controlUnit;

ARCHITECTURE Behavioral OF controlUnit IS
    TYPE procStateType IS (SETUP, FETCH_SETUP, FETCH_MEM_READ, DECODE, EXECUTE, MEM_ACCESS, WRITE_BACK);
    SIGNAL procState, procState_nxt : procStateType;

    --internal registers
    SIGNAL currentlyHandlingInterruptReg, currentlyHandlingInterruptReg_nxt           : BOOLEAN;
    SIGNAL currentlyHandlingInterruptIndexReg, currentlyHandlingInterruptIndexReg_nxt : unsigned(7 DOWNTO 0);
    SIGNAL currentInterruptHandlerAddressReg, currentInterruptHandlerAddressReg_nxt   : STD_LOGIC_VECTOR(31 DOWNTO 0);

    SIGNAL currentlyHaltingReg, currentlyHaltingReg_nxt : BOOLEAN;

    SIGNAL softwareResetReg, softwareResetReg_nxt : STD_LOGIC := '0';

    --signals to keep track of decoded information within instructions
    SIGNAL instructionReg, instructionReg_nxt                             : STD_LOGIC_VECTOR(31 DOWNTO 0);
    SIGNAL destinationRegisterNumberReg, destinationRegisterNumberReg_nxt : INTEGER;
    SIGNAL addressRegisterNumberReg, addressRegisterNumberReg_nxt         : INTEGER;
    SIGNAL sourceRegisterNumberReg, sourceRegisterNumberReg_nxt           : INTEGER;
    SIGNAL useCPSR_EnReg, useCPSR_EnReg_nxt                               : BOOLEAN;
    SIGNAL writeBackEnReg, writeBackEnReg_nxt                             : BOOLEAN;
    SIGNAL writeFromALU_EnReg, writeFromALU_EnReg_nxt                     : BOOLEAN;
    SIGNAL updateCPSR_EnReg, updateCPSR_EnReg_nxt                         : BOOLEAN;
    SIGNAL writeAddressBackEnReg, writeAddressBackEnReg_nxt               : BOOLEAN;
    SIGNAL memOperationReg, memOperationReg_nxt                           : STD_LOGIC; --1: read, 0: write

    SIGNAL CPSR_Reg, CPSR_Reg_nxt           : STD_LOGIC_VECTOR(3 DOWNTO 0);
    SIGNAL CPSR_Reg_Temp, CPSR_Reg_Temp_nxt : STD_LOGIC_VECTOR(3 DOWNTO 0);
    SIGNAL PC_Reg_Temp, PC_Reg_Temp_nxt     : STD_LOGIC_VECTOR(31 DOWNTO 0);

    SIGNAL Z_flag : STD_LOGIC;
    SIGNAL N_flag : STD_LOGIC;
    SIGNAL V_flag : STD_LOGIC;
    SIGNAL C_flag : STD_LOGIC;

    --registers that keep track of the control signals of the ALU (only the control Signal for the ALU need a separate register) 
    SIGNAL operand1SelReg, operand1SelReg_nxt                     : STD_LOGIC_VECTOR(4 DOWNTO 0) := (OTHERS => '0');
    SIGNAL operand2SelReg, operand2SelReg_nxt                     : STD_LOGIC_VECTOR(4 DOWNTO 0) := (OTHERS => '0');
    SIGNAL bitManipulationValSelReg, bitManipulationValSelReg_nxt : STD_LOGIC_VECTOR(4 DOWNTO 0) := (OTHERS => '0');
    SIGNAL bitManipulationCodeReg, bitManipulationCodeReg_nxt     : STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
    SIGNAL bitManipulationValueReg, bitManipulationValueReg_nxt   : STD_LOGIC_VECTOR(4 DOWNTO 0) := (OTHERS => '0');

    SIGNAL ALU_opCodeReg, ALU_opCodeReg_nxt : STD_LOGIC_VECTOR(3 DOWNTO 0)  := (OTHERS => '0');
    SIGNAL carryInReg, carryInReg_nxt       : STD_LOGIC                     := '0';
    SIGNAL upperSelReg, upperSelReg_nxt     : STD_LOGIC                     := '0';
    SIGNAL dataToALU_Reg, dataToALU_Reg_nxt : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');

    --delay register
    SIGNAL delayReg, delayReg_nxt : STD_LOGIC;

    --interrupt registers
    SIGNAL invalidInstructionInterruptReg, invalidInstructionInterruptReg_nxt : STD_LOGIC;
    SIGNAL softwareInterruptReg, softwareInterruptReg_nxt                     : STD_LOGIC;

    --bit masks
    TYPE bitMasksType IS ARRAY (0 TO 16) OF STD_LOGIC_VECTOR(31 DOWNTO 0);

    CONSTANT bitMasks : bitMasksType := (
        0  => x"00000000",
        1  => x"00000001",
        2  => x"00000003",
        3  => x"0000000F",
        4  => x"000000FF",
        5  => x"0000FF00",
        6  => x"0F0F0F0F",
        7  => x"F0F0F0F0",
        8  => x"55555555",
        9  => x"AAAAAAAA",
        10 => x"FFFFFFFF",
        OTHERS => (OTHERS => '0')
    );

    --operation codes
    --Data Processing
    CONSTANT ANDD : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
    CONSTANT EOR  : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0001";
    CONSTANT ORR  : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0010";
    CONSTANT BIC  : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0011";
    CONSTANT NOTT : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0100";
    CONSTANT SUB  : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0101";
    CONSTANT BUSS : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0110";
    CONSTANT ADDD : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0111";
    CONSTANT ADC  : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1000";
    CONSTANT SBC  : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1001";
    CONSTANT BSC  : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1010";
    CONSTANT MOV  : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1011";
    CONSTANT MUL  : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1100";
    CONSTANT UMUL : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1101";

    --Data Movement 
    CONSTANT LOAD  : STD_LOGIC_VECTOR(2 DOWNTO 0) := "000";
    CONSTANT STORE : STD_LOGIC_VECTOR(2 DOWNTO 0) := "001";

    --Special Instructions
    CONSTANT PASS : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
    CONSTANT HALT : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0001";
    CONSTANT SIR  : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0010";
    CONSTANT RES  : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0011";
    CONSTANT IRET : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0100";

    CONSTANT IINIT : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1111"; --this is an internal instruction that initializes an interrupt handler. It cannot be used in assembly language.
    --Control Flow 
    CONSTANT JUMP  : STD_LOGIC_VECTOR(1 DOWNTO 0) := "00";
    CONSTANT JUMPL : STD_LOGIC_VECTOR(1 DOWNTO 0) := "01";

    --Booloader code. This code is executed when programming mode is enabled.
    TYPE ROM IS ARRAY (0 TO 256) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
    CONSTANT bootloaderMemory : ROM := (
        0  => "11111101110000000000101000001011",
        1  => "11111101111010000000000000001100",
        2  => "11111001000000000000110010111011",
        3  => "11111101110001001000011010001010",
        4  => "11111101111000000001111010001100",
        5  => "11111001000000000000110010101010",
        6  => "11110000100000000000000010111010",
        7  => "11111101110000000000000000000000",
        8  => "11110110110000000000000000011010",
        9  => "11111101110000000000110000001010",
        10 => "11111101111010000000000000001100",
        11 => "11111001000000000000110010101010",
        12 => "11110000000000000000000010101001",
        13 => "11111101100100001000000100101001",
        14 => "11111010111000000000100101000000",
        15 => "00010110011000000000000000000111",
        16 => "11111101110000000000000000000001",
        17 => "11111101110000000000000000000010",
        18 => "11111101110000000000110010001010",
        19 => "11111101111010000000000000001100",
        20 => "11111001000000000000110010101010",
        21 => "11110000000000000000000010101001",
        22 => "11111101110000000010000000001010",
        23 => "11111000001000000000100110100000",
        24 => "00010110010000000000000000010100",
        25 => "11111101100010000110000000100011",
        26 => "11111001000011000110001010010010",
        27 => "11111011110000000000000100010001",
        28 => "11111010111000000000000101000000",
        29 => "00010110011000000000000000001100",
        30 => "11110000100000000000000000000010",
        31 => "11111011110000000000000001000000",
        32 => "11111101110000000001111111101000",
        33 => "11110110110000000000000000000110",
        34 => "11110110011000000000000000011011",
        35 => "11111101110000000000101010000110",
        36 => "11111101111010000000000000001100",
        37 => "11111001000000000000110001100110",
        38 => "11110000100000000000000001100000",
        39 => "11111101100000000000000110101111",
        40 => "11111101110000000000110010000110",
        41 => "11111101111010000000000000001100",
        42 => "11111001000000000000110001100110",
        43 => "11110000100000000000000001101000",
        44 => "11111101100000000000000110101111",
        45 => "11111101110000000001000000001000",
        46 => "11110110111000000000000000000111",
        47 => "11110110011000000000000000101000",
        OTHERS => (OTHERS => '0')
    );

BEGIN
    --assigning interrupt signals
    interrupts(0) <= invalidInstructionInterruptReg;
    interrupts(1) <= softwareInterruptReg;

    --assigning debug signals
    debug(38 DOWNTO 7) <= instructionReg;
    debug(6)           <= Z_flag;
    debug(5)           <= N_flag;
    debug(4)           <= V_flag;
    debug(3)           <= C_flag;

    convertingStateToDebugSignal : PROCESS (procState)
        VARIABLE bitRepresentationState : STD_LOGIC_VECTOR(2 DOWNTO 0);
    BEGIN
        CASE procState IS
            WHEN SETUP          => bitRepresentationState          := "000";
            WHEN FETCH_SETUP    => bitRepresentationState    := "001";
            WHEN FETCH_MEM_READ => bitRepresentationState := "010";
            WHEN DECODE         => bitRepresentationState         := "011";
            WHEN EXECUTE        => bitRepresentationState        := "100";
            WHEN MEM_ACCESS     => bitRepresentationState     := "101";
            WHEN WRITE_BACK     => bitRepresentationState     := "110";
            WHEN OTHERS         => bitRepresentationState         := "000";
        END CASE;
        debug(2 DOWNTO 0) <= bitRepresentationState;
    END PROCESS;

    --assigning flag signals
    Z_flag <= CPSR_Reg(3);
    N_flag <= CPSR_Reg(2);
    V_flag <= CPSR_Reg(1);
    C_flag <= CPSR_Reg(0);

    stateMachine : PROCESS (PC, procState, interruptIndex, currentInterruptHandlerAddressReg, PC_Reg_Temp, CPSR_Reg_Temp, currentlyHandlingInterruptIndexReg, operand1SelReg, operand2SelReg, bitManipulationValSelReg, bitManipulationCodeReg, bitManipulationValueReg, ALU_opCodeReg, carryInReg, upperSelReg, dataToALU_Reg, programmingMode, InterruptHandlerAddress, dataFromMem, dataFromALU, flagsFromALU, memOpFinished, instructionReg, destinationRegisterNumberReg, useCPSR_EnReg, writeBackEnReg, writeFromALU_EnReg, updateCPSR_EnReg, memOperationReg, addressRegisterNumberReg, writeAddressBackEnReg, sourceRegisterNumberReg, CPSR_Reg, Z_flag, N_flag, V_flag, C_flag, softwareInterruptReg, invalidInstructionInterruptReg, currentlyHandlingInterruptReg, currentlyHaltingReg, delayReg, softwareResetReg)
        VARIABLE condition    : STD_LOGIC_VECTOR(3 DOWNTO 0);
        VARIABLE conditionMet : STD_LOGIC;
        TYPE instructionClassType IS (DATA_PROCESSING, DATA_MOVEMENT, SPECIAL, CONTROL_FLOW, INVALID);
        VARIABLE instructionClass : instructionClassType;

        --variables for the different instruction classes:
        --Data Processing
        VARIABLE dataProcessingInstructionOpCode : STD_LOGIC_VECTOR(3 DOWNTO 0);

        --Data Movement
        VARIABLE dataMovementInstructionOpCode : STD_LOGIC_VECTOR(2 DOWNTO 0);

        --Special Instructions
        VARIABLE specialInstructionOpCode : STD_LOGIC_VECTOR(3 DOWNTO 0);

        --Control Flow
        VARIABLE controlFlowInstructionOpCode : STD_LOGIC_VECTOR(1 DOWNTO 0);

        --variables for different sections within the instruction:
        VARIABLE sourceReg       : STD_LOGIC_VECTOR(3 DOWNTO 0);
        VARIABLE addressRegister : STD_LOGIC_VECTOR(3 DOWNTO 0);
        VARIABLE immediateEn     : STD_LOGIC;
        VARIABLE offsetEn        : STD_LOGIC;
        VARIABLE offset          : STD_LOGIC_VECTOR(11 DOWNTO 0);
        VARIABLE subtractEn      : STD_LOGIC;
        VARIABLE immediateValue  : STD_LOGIC_VECTOR(31 DOWNTO 0);

        VARIABLE bitManipulationMethod   : STD_LOGIC_VECTOR(1 DOWNTO 0);
        VARIABLE bitManipulationUseRegEn : STD_LOGIC;
        VARIABLE bitManipulationOperand  : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
        --default assignments for control signals
        operand1Sel           <= (OTHERS => '1');
        operand2Sel           <= (OTHERS => '1');
        dataToMemSel          <= (OTHERS => '0');
        dataToRegistersSel    <= '0';
        bitManipulationValSel <= (OTHERS => '1');
        loadRegistersSel      <= (OTHERS => '0');
        interruptsClr         <= (OTHERS => '0');
        bitManipulationCode   <= (OTHERS => '0');
        bitManipulationValue  <= (OTHERS => '0');
        ALU_opCode            <= (OTHERS => '0');
        carryIn               <= '0';
        upperSel              <= '0';
        memWriteReq           <= '0';
        memReadReq            <= '0';
        dataToALU             <= (OTHERS => '0');
        ALU_En                <= '0';
        createLink            <= '0';

        --controlRegisters
        instructionReg_nxt                     <= instructionReg;
        procState_nxt                          <= procState;
        CPSR_Reg_nxt                           <= CPSR_Reg;
        CPSR_Reg_Temp_nxt                      <= CPSR_Reg_Temp;
        PC_Reg_Temp_nxt                        <= PC_Reg_Temp;
        invalidInstructionInterruptReg_nxt     <= invalidInstructionInterruptReg;
        softwareInterruptReg_nxt               <= softwareInterruptReg;
        currentlyHandlingInterruptReg_nxt      <= currentlyHandlingInterruptReg;
        currentlyHandlingInterruptIndexReg_nxt <= currentlyHandlingInterruptIndexReg;
        currentInterruptHandlerAddressReg_nxt  <= currentInterruptHandlerAddressReg;
        currentlyHaltingReg_nxt                <= currentlyHaltingReg;

        --temporary registers for holding information about the current instruction
        destinationRegisterNumberReg_nxt <= destinationRegisterNumberReg;
        addressRegisterNumberReg_nxt     <= addressRegisterNumberReg;
        useCPSR_EnReg_nxt                <= useCPSR_EnReg;
        writeBackEnReg_nxt               <= writeBackEnReg;
        writeFromALU_EnReg_nxt           <= writeFromALU_EnReg;
        updateCPSR_EnReg_nxt             <= updateCPSR_EnReg;
        memOperationReg_nxt              <= memOperationReg;
        writeAddressBackEnReg_nxt        <= writeAddressBackEnReg;
        sourceRegisterNumberReg_nxt      <= sourceRegisterNumberReg;

        --registers that save the state of the control signals of the ALU
        operand1SelReg_nxt           <= operand1SelReg;
        operand2SelReg_nxt           <= operand2SelReg;
        bitManipulationValSelReg_nxt <= bitManipulationValSelReg;
        bitManipulationCodeReg_nxt   <= bitManipulationCodeReg;
        bitManipulationValueReg_nxt  <= bitManipulationValueReg;
        ALU_opCodeReg_nxt            <= ALU_opCodeReg;
        carryInReg_nxt               <= carryInReg;
        upperSelReg_nxt              <= upperSelReg;
        dataToALU_Reg_nxt            <= dataToALU_Reg;

        --delay register
        delayReg_nxt <= delayReg;

        --reset register
        softwareResetReg_nxt <= softwareResetReg;

        IF procState = SETUP THEN
            procState_nxt <= FETCH_SETUP;
            --set ALU signal registers for the next instruction fetch
            operand2SelReg_nxt <= "01111"; --selecting PC as operand 2
            ALU_opCodeReg_nxt  <= "1011";  --tell ALU to MOV PC to output.

        ELSIF procState = FETCH_SETUP THEN
            IF NOT(unsigned(interruptHandlerAddress) /= 0 AND currentlyHandlingInterruptReg = False) THEN
                IF currentlyHaltingReg = False THEN
                    procState_nxt <= FETCH_MEM_READ;

                    --set ALU control signals
                    operand2Sel <= operand2SelReg;
                    ALU_opCode  <= ALU_opCodeReg;

                    --enable ALU
                    ALU_En <= '1';

                    --Prepare ALU control signals for next state, where the PC will be incremented.
                    operand1SelReg_nxt <= "10000";     --dataToALU as operand 1.
                    operand2SelReg_nxt <= "01111";     --Selecting PC as operand 2.
                    dataToALU_Reg_nxt  <= x"00000004"; --set dataToALU to 4 to increment PC later
                    ALU_opCodeReg_nxt  <= "0111";      --tell ALU to add operand1 (4) to the PC
                ELSE
                    procState_nxt <= FETCH_SETUP;
                END IF;

            ELSE
                --an interrupt has occured and the interrupt handler will now be initialized.
                currentlyHaltingReg_nxt                <= False;
                currentlyHandlingInterruptReg_nxt      <= True;
                instructionReg_nxt                     <= "11110101111000000000000000000000";
                currentInterruptHandlerAddressReg_nxt  <= interruptHandlerAddress;
                currentlyHandlingInterruptIndexReg_nxt <= unsigned(interruptIndex);
                procState_nxt                          <= DECODE;

            END IF;

        ELSIF procState = FETCH_MEM_READ THEN
            memReadReq  <= '1';
            operand1Sel <= operand1SelReg;
            operand2Sel <= operand2SelReg;
            dataToALU   <= dataToALU_Reg;
            ALU_opCode  <= ALU_opCodeReg;
            --Handle instruction fetch in programming mode.
            IF programmingMode = '1' THEN
                instructionReg_nxt <= bootloaderMemory(to_integer(unsigned(dataFromALU(9 DOWNTO 2)))); --Address needs to be divided by four.
                ALU_En             <= '1';                                                             --enable ALU in order to increment the PC
                procState_nxt      <= DECODE;

                --Handle instruction fetch in normal mode.
            ELSE
                IF memOpFinished = '1' THEN        --wait for data to arrive         
                    instructionReg_nxt <= dataFromMem; --load current instruction into the instruction register
                    ALU_En             <= '1';         --enable ALU in order to increment the PC
                    procState_nxt      <= DECODE;
                END IF;
            END IF;
        ELSIF procState = DECODE THEN
            loadRegistersSel   <= "1000000000000000"; --load value back into PC
            dataToRegistersSel <= '0';                --sending data from ALU to registers in order to write the incremented address back to the PC

            procState_nxt <= EXECUTE; --The next state will always be "EXECUTE" state.

            --default assignments
            operand1SelReg_nxt           <= (OTHERS => '0');
            operand2SelReg_nxt           <= (OTHERS => '0');
            bitManipulationValSelReg_nxt <= (OTHERS => '1');
            bitManipulationCodeReg_nxt   <= (OTHERS => '0');
            bitManipulationValueReg_nxt  <= (OTHERS => '0');
            ALU_opCodeReg_nxt            <= (OTHERS => '0');
            carryInReg_nxt               <= '0'; --not used yet
            upperSelReg_nxt              <= '0'; --not used yet
            dataToALU_Reg_nxt            <= (OTHERS => '0');

            --extract condition from instruction
            condition := instructionReg(31 DOWNTO 28);
            CASE condition IS
                WHEN "0000" => conditionMet := Z_flag;                                  --equal
                WHEN "0001" => conditionMet := NOT Z_flag;                              --not equal
                WHEN "0010" => conditionMet := C_flag;                                  --unsigned higher or same
                WHEN "0011" => conditionMet := NOT C_flag;                              --unsigned lower
                WHEN "0100" => conditionMet := N_flag;                                  --negative
                WHEN "0101" => conditionMet := NOT N_flag;                              --positive or zero
                WHEN "0110" => conditionMet := V_flag;                                  --overflow
                WHEN "0111" => conditionMet := NOT V_flag;                              --no overflow
                WHEN "1000" => conditionMet := C_flag AND (NOT Z_flag);                 -- unsigned higher
                WHEN "1001" => conditionMet := (NOT C_flag) OR Z_flag;                  --unsigned lower or same
                WHEN "1010" => conditionMet := NOT (N_flag XOR V_flag);                 --greater or equal
                WHEN "1011" => conditionMet := N_flag XOR V_flag;                       --less than
                WHEN "1100" => conditionMet := (NOT Z_flag) AND NOT(N_flag XOR V_flag); --greater than
                WHEN "1101" => conditionMet := (NOT Z_flag) OR (N_flag XOR V_flag);     --less than or equal
                WHEN OTHERS => conditionMet := '1';                                     --always
            END CASE;

            --skip instruction if condition is not met
            IF NOT conditionMet = '1' THEN
                --set ALU signal registers for the next instruction fetch
                operand2SelReg_nxt <= "01111"; --selecting PC as operand 2
                ALU_opCodeReg_nxt  <= "1011";  --tell ALU to MOV PC to output.
                procState_nxt      <= FETCH_SETUP;
            ELSE
                --IF an instruction uses bit manipulation, it will ALWAYS use bit 20-13. Therefore, it can be set in the beginning without any conditions. However, each instruction sets "bitManipulationValSel" individually depending on whether (and if yes how) it  uses bit manipulation. Setting "bitManipulationValSel="11111"" will tell the ALU to not make use of bit manipulation.
                bitManipulationMethod   := instructionReg(20 DOWNTO 19);
                bitManipulationUseRegEn := instructionReg(18);
                bitManipulationOperand  := instructionReg(17 DOWNTO 13);
                bitManipulationCodeReg_nxt  <= bitManipulationMethod;
                bitManipulationValueReg_nxt <= bitManipulationOperand;

                --check what kind of instruction class the instruction belongs to
                IF instructionReg(27) = '1' THEN
                    instructionClass := DATA_PROCESSING;
                ELSIF instructionReg(27 DOWNTO 26) = "00" THEN
                    instructionClass := DATA_MOVEMENT;
                ELSIF instructionReg(27 DOWNTO 25) = "010" THEN
                    instructionClass := SPECIAL;
                ELSIF instructionReg(27 DOWNTO 25) = "011" THEN
                    instructionClass := CONTROL_FLOW;
                ELSE
                    instructionClass := INVALID;               --needs to be set to avoid latch
                    invalidInstructionInterruptReg_nxt <= '1'; --handle invalid instructions
                    procState_nxt                      <= SETUP;
                END IF;
                --handle different instructin classes 
                CASE instructionClass IS
                    WHEN DATA_PROCESSING =>
                        updateCPSR_EnReg_nxt   <= True;--All of the Data Processing instructions (except MOV) update the CPSR register.
                        useCPSR_EnReg_nxt      <= False; --this is a default assignments, in some cases the CPSR will be used as the destination register.
                        writeBackEnReg_nxt     <= True;  --This instruction class always writes back to register file.
                        writeFromALU_EnReg_nxt <= True;  --This instruction class updates registers from ALU result.

                        destinationRegisterNumberReg_nxt <= to_integer(unsigned(instructionReg(3 DOWNTO 0))); --All instructions in this instruction class use the same bits for the destination Register.

                        immediateEn := instructionReg(22);--All instructions in this instruction class use the same bit as their "Immediate Enable Bit".

                        dataProcessingInstructionOpCode := instructionReg(26 DOWNTO 23);
                        ALU_opCodeReg_nxt <= dataProcessingInstructionOpCode; --Tell ALU which operation to perform.

                        IF dataProcessingInstructionOpCode = MOV THEN --the MOV instruction is different from the other ones.
                            updateCPSR_EnReg_nxt <= False;
                            IF instructionReg(4) = '1' THEN --if this bit is set, the destination register is the CPSR.
                                useCPSR_EnReg_nxt <= True;
                            END IF;

                            IF immediateEn = '1' THEN
                                IF instructionReg(21) = '1' THEN --checks if the "Load Higher Bytes Enable Bit" is set.
                                    immediateValue := instructionReg(20 DOWNTO 5) & x"0000";
                                ELSE
                                    immediateValue := x"0000" & instructionReg(20 DOWNTO 5);
                                END IF;
                                operand2SelReg_nxt <= "10000"; --tells the ALU to use "dataToALU" as operand 2.
                                dataToALU_Reg_nxt  <= immediateValue;
                            ELSE
                                operand2SelReg_nxt <= instructionReg(9 DOWNTO 5);
                                IF instructionReg(9) = '1' THEN --if this bit is set, the source register is the CPSR.
                                    dataToALU_Reg_nxt <= x"0000000" & CPSR_Reg;
                                END IF;
                                IF bitManipulationUseRegEn = '0' THEN
                                    bitManipulationValSelReg_nxt <= "10000"; --uses the "bitManipulationOperand" as immediate value for bit manipulation.
                                ELSE
                                    bitManipulationValSelReg_nxt <= '0' & bitManipulationOperand(3 DOWNTO 0); --uses the "bitManipulationOperand" as register for bit manipulation
                                END IF;

                            END IF;
                        ELSE
                            --all of these instruction will always apply bit manipulation to operand 2
                            IF bitManipulationUseRegEn = '0' THEN
                                bitManipulationValSelReg_nxt <= "10000"; --uses the "bitManipulationOperand" as immediate value for bit manipulation.
                            ELSE
                                bitManipulationValSelReg_nxt <= '0' & bitManipulationOperand(3 DOWNTO 0); --uses the "bitManipulationOperand" as register for bit manipulation
                            END IF;

                            --all instruction specify the operand 1 register in the same way
                            operand1SelReg_nxt <= '0' & instructionReg(11 DOWNTO 8);

                            --all instructions use the same bit to tell the cpu, if operand 2 should be interpreted as a register or as something else.      
                            IF immediateEn = '1' THEN
                                operand2SelReg_nxt <= "10000"; --operand 2 will be specified by CU
                            ELSE
                                operand2SelReg_nxt <= '0' & instructionReg(7 DOWNTO 4); --operand 2 will be a register
                            END IF;
                            IF dataProcessingInstructionOpCode = ANDD OR dataProcessingInstructionOpCode = EOR OR dataProcessingInstructionOpCode = ORR OR dataProcessingInstructionOpCode = BIC OR dataProcessingInstructionOpCode = NOTT THEN
                                --These instructions do not offer the possibility to specify immediate values. Instead, a bit mask can be specified.
                                IF immediateEn = '1' THEN
                                    dataToALU_Reg_nxt <= bitMasks(to_integer(unsigned(instructionReg(7 DOWNTO 4))));
                                END IF;
                                --These instructions can disable write back if bit 21 of the instruction is set.
                                IF instructionReg(21) = '1' THEN
                                    writeBackEnReg_nxt <= False;
                                END IF;

                            ELSIF dataProcessingInstructionOpCode = SUB OR dataProcessingInstructionOpCode = BUSS OR dataProcessingInstructionOpCode = ADDD OR dataProcessingInstructionOpCode = ADC OR dataProcessingInstructionOpCode = SBC OR dataProcessingInstructionOpCode = BSC THEN
                                --These instructions offer you to specify an immediate value.
                                IF immediateEn = '1' THEN
                                    dataToALU_Reg_nxt <= x"0000000" & instructionReg(7 DOWNTO 4);
                                END IF;

                                --These instructions can disable write back if bit 21 of the instruction is set.
                                IF instructionReg(21) = '1' THEN
                                    writeBackEnReg_nxt <= False;
                                END IF;

                            ELSIF dataProcessingInstructionOpCode = MUL OR dataProcessingInstructionOpCode = UMUL THEN
                                --These instructions offer you to specify an immediate value.
                                IF immediateEn = '1' THEN
                                    dataToALU_Reg_nxt <= x"0000000" & instructionReg(7 DOWNTO 4);
                                END IF;
                                --Since these instructions perform multiplications, it needs to be specified, whether to write back the upper or lower 32 bits of the result.
                                upperSelReg_nxt <= instructionReg(21);
                            ELSE
                                invalidInstructionInterruptReg_nxt <= '1';
                            END IF;

                        END IF;
                    WHEN DATA_MOVEMENT =>
                        dataMovementInstructionOpCode := instructionReg(25 DOWNTO 23);
                        updateCPSR_EnReg_nxt      <= False;--None of the Data Processing instructions update the CPSR register.
                        useCPSR_EnReg_nxt         <= False; --None of the Data Movement instructions update the status flags.
                        writeBackEnReg_nxt        <= True;  --This instruction class always updates the registers.
                        writeFromALU_EnReg_nxt    <= False; --This instruction class updates registers from memory.
                        writeAddressBackEnReg_nxt <= False; --This is a default assignment. In some cases the altered address will be written back to the addressRegister.

                        IF dataMovementInstructionOpCode = STORE OR dataMovementInstructionOpCode = LOAD THEN
                            --differentiate between load and store instruction
                            IF dataMovementInstructionOpCode = STORE THEN
                                memOperationReg_nxt         <= '0';
                                sourceRegisterNumberReg_nxt <= to_integer(unsigned(instructionReg(3 DOWNTO 0))); --CAN BE REMOVED???
                            ELSE
                                memOperationReg_nxt              <= '1';
                                destinationRegisterNumberReg_nxt <= to_integer(unsigned(instructionReg(3 DOWNTO 0)));
                            END IF;

                            --otherwise, the two instructions work exactly the same:
                            addressRegister := instructionReg(7 DOWNTO 4);
                            addressRegisterNumberReg_nxt <= to_integer(unsigned(addressRegister));
                            operand2SelReg_nxt           <= '0' & addressRegister; --operand 2 will be data in specified register.
                            operand1SelReg_nxt           <= "10000";               --operand one will be the data sent by control unit.

                            offsetEn := instructionReg(21);
                            IF offsetEn = '1' THEN
                                subtractEn := instructionReg(20);
                                offset     := instructionReg(19 DOWNTO 8);
                                dataToALU_Reg_nxt <= x"00000" & offset;
                                --subtract or add the offset to the current
                                IF subtractEn = '1' THEN
                                    ALU_opCodeReg_nxt <= "0110"; --operation code for subraction (operand2 - operand1)
                                ELSE
                                    ALU_opCodeReg_nxt <= "0111"; --operation code for addition (operand2 + operand 1)
                                END IF;
                            ELSE
                                --ignore operand 1
                                ALU_opCodeReg_nxt <= "1011";
                                --Apply bit manipulation to operand2.
                                IF bitManipulationUseRegEn = '0' THEN
                                    bitManipulationValSelReg_nxt <= "10000"; --Uses the "bitManipulationOperand" as immediate value for bit manipulation.
                                ELSE
                                    bitManipulationValSelReg_nxt <= '0' & bitManipulationOperand(3 DOWNTO 0); --uses the "bitManipulationOperand" as register for bit manipulation.
                                END IF;
                            END IF;
                            IF instructionReg(22) = '1' THEN
                                writeAddressBackEnReg_nxt <= True;
                            END IF;
                        ELSE
                            invalidInstructionInterruptReg_nxt <= '1'; --handle invalid instructions
                            procState_nxt                      <= SETUP;
                        END IF;

                    WHEN SPECIAL =>
                        specialInstructionOpCode := instructionReg(24 DOWNTO 21);
                        --default assignments
                        updateCPSR_EnReg_nxt <= False;--None of the Data Processing instructions update the CPSR register.
                        useCPSR_EnReg_nxt    <= False; --None of the Data Movement instructions update the status flags.
                        writeBackEnReg_nxt   <= False; --Only the Interrupt Init Instruction needs a register write back.

                        --Set ALU signal registers for the next instruction fetch for those instructions that dont need memeory access and write back.
                        operand2SelReg_nxt <= "01111"; --Selecting PC as operand 2
                        ALU_opCodeReg_nxt  <= "1011";  --Tell ALU to MOV PC to output.
                        procState_nxt      <= FETCH_SETUP;

                        --check if the remaining Bits are zero
                        IF instructionReg(20 DOWNTO 0) = "000000000000000000000" THEN
                            CASE specialInstructionOpCode IS
                                WHEN PASS =>
                                    NULL;
                                WHEN HALT =>
                                    currentlyHaltingReg_nxt <= True;

                                WHEN SIR =>
                                    softwareInterruptReg_nxt <= '1';

                                WHEN IRET =>
                                    currentlyHandlingInterruptReg_nxt <= False;
                                    CPSR_Reg_nxt                      <= CPSR_Reg_Temp; --Restore flags.

                                    --Prepare Restoring PC.
                                    operand2SelReg_nxt               <= "10000";
                                    dataToALU_Reg_nxt                <= PC_Reg_Temp;
                                    writeBackEnReg_nxt               <= True;
                                    writeFromALU_EnReg_nxt           <= True;
                                    destinationRegisterNumberReg_nxt <= 15;
                                    procState_nxt                    <= EXECUTE;

                                WHEN IINIT =>
                                    --Clear The interrupt at the beginning of the interrupt handler routine. 
                                    IF currentlyHandlingInterruptIndexReg = 0 THEN
                                        invalidInstructionInterruptReg_nxt <= '0';
                                    ELSIF currentlyHandlingInterruptIndexReg = 1 THEN
                                        softwareInterruptReg_nxt <= '0';
                                    ELSIF currentlyHandlingInterruptIndexReg < numInterrupts THEN
                                        interruptsClr(to_integer(currentlyHandlingInterruptIndexReg) - 2) <= '1';
                                    ELSE
                                        NULL;
                                    END IF;

                                    CPSR_Reg_Temp_nxt                <= CPSR_Reg; --Save current flags                
                                    PC_Reg_Temp_nxt                  <= PC;       --Save current PC
                                    operand2SelReg_nxt               <= "10000";  --tells the ALU to use "dataToALU" as operand 2.
                                    dataToALU_Reg_nxt                <= currentInterruptHandlerAddressReg;
                                    writeBackEnReg_nxt               <= True;
                                    writeFromALU_EnReg_nxt           <= True;
                                    destinationRegisterNumberReg_nxt <= 15; --Write Result into PC
                                    procState_nxt                    <= EXECUTE;

                                WHEN RES =>
                                    softwareResetReg_nxt <= '1';

                                WHEN OTHERS =>
                                    invalidInstructionInterruptReg_nxt <= '1'; --Handle invalid instructions.
                            END CASE;
                        ELSE
                            invalidInstructionInterruptReg_nxt <= '1'; --Handle invalid instructions.
                        END IF;

                    WHEN CONTROL_FLOW =>
                        controlFlowInstructionOpCode := instructionReg(24 DOWNTO 23);
                        updateCPSR_EnReg_nxt   <= False;--None of the Data Processing instructions update the CPSR register.
                        useCPSR_EnReg_nxt      <= False; --The CPSR Register cannnot be used as a parameter. 
                        writeBackEnReg_nxt     <= True;  --This instruction class always updates the registers.
                        writeFromALU_EnReg_nxt <= True;  --This instruction class updates registers from the ALU.
                        IF controlFlowInstructionOpCode = JUMP OR controlFlowInstructionOpCode = JUMPL THEN
                            --The program counter is always the source register 
                            destinationRegisterNumberReg_nxt <= 15;
                            createLink                       <= controlFlowInstructionOpCode(0); --Only create a link if the op code belongs to the JUMPL instruction.

                            --set the ALU signals
                            operand1SelReg_nxt <= "01111";                                          --Select PC as operand 1.
                            IF instructionReg(22) = '1' THEN                                        --Check if 'Immediate Offset Enable Bit' is set.
                                operand2SelReg_nxt <= "10000";                                          --Select data from CU as operand 2.
                                dataToALU_Reg_nxt  <= "000000000" & instructionReg(20 DOWNTO 0) & "00"; --Multiply immediate value by 4 (so that it is a valid memory address) and send it to ALU.
                                IF instructionReg(21) = '1' THEN                                        --Check if the 'Subtract Bit' is set.
                                    ALU_opCodeReg_nxt <= "0101";                                            --ALU operation Code for subtraction.
                                ELSE
                                    ALU_opCodeReg_nxt <= "0111"; --ALU operation Code for addition.
                                END IF;
                            ELSE
                                operand2SelReg_nxt <= '0' & instructionReg(3 DOWNTO 0); --Select specified register as operand 2.
                                IF bitManipulationUseRegEn = '0' THEN
                                    bitManipulationValSelReg_nxt <= "10000"; --uses the "bitManipulationOperand" as immediate value for bit manipulation.
                                ELSE
                                    bitManipulationValSelReg_nxt <= '0' & bitManipulationOperand(3 DOWNTO 0); --uses the "bitManipulationOperand" as register for bit manipulation
                                END IF;
                                IF instructionReg(21) = '1' THEN --Check if the 'Register as Offset Enable Bit' is set.
                                    ALU_opCodeReg_nxt <= "0111";     --ALU operation Code for addition (offset will be added to the PC)
                                ELSE
                                    ALU_opCodeReg_nxt <= "1011"; --ALU operation Code for MOV (The value of operand2 will be copied into the PC).
                                END IF;
                            END IF;
                        ELSE
                            invalidInstructionInterruptReg_nxt <= '1'; --Handle invalid instructions.
                        END IF;

                    WHEN OTHERS =>
                        invalidInstructionInterruptReg_nxt <= '1'; --Handle invalid instructions.
                        procState_nxt                      <= SETUP;
                END CASE;
            END IF;

        ELSIF procState = Execute THEN
            ALU_En                <= '1'; --enable ALU
            operand1Sel           <= operand1SelReg;
            operand2Sel           <= operand2SelReg;
            bitManipulationValSel <= bitManipulationValSelReg;
            bitManipulationCode   <= bitManipulationCodeReg;
            bitManipulationValue  <= bitManipulationValueReg;
            ALU_opCode            <= ALU_opCodeReg;
            carryIn               <= carryInReg;
            upperSel              <= upperSelReg;
            dataToALU             <= dataToALU_Reg;

            --wait one clock cycle for the result and the flags to arrive
            IF delayReg = '1' THEN
                IF writeFromALU_EnReg = True THEN
                    procState_nxt <= WRITE_BACK;
                ELSE
                    procState_nxt <= MEM_ACCESS;
                END IF;
                delayReg_nxt <= '0';
            ELSE
                delayReg_nxt <= '1';
            END IF;
        ELSIF procState = MEM_ACCESS THEN
            IF memOperationReg = '1' THEN --read
                memReadReq    <= '1';
                procState_nxt <= WRITE_BACK; --After loading a value from memory, that value needs to be written to a register. 
            ELSE
                memWriteReq <= '1'; --write
                IF memOpFinished = '1' THEN
                    procState_nxt <= FETCH_SETUP; --After storing a value in memory, No register access will be needed.
                END IF;
            END IF;
            dataToMemSel <= STD_LOGIC_VECTOR(to_unsigned(sourceRegisterNumberReg, 4));

            IF writeAddressBackEnReg = True THEN
                loadRegistersSel(addressRegisterNumberReg) <= '1'; --Select address register as write back register.
                dataToRegistersSel                         <= '0'; --Load registers from ALU output.
            END IF;

            --set ALU signal registers for the next instruction fetch
            operand2SelReg_nxt <= "01111"; --selecting PC as operand 2
            ALU_opCodeReg_nxt  <= "1011";  --tell ALU to MOV PC to output.

        ELSIF procState = WRITE_BACK THEN
            --default assignment
            procState_nxt <= FETCH_SETUP;

            --Handling the updates of the status flags.
            IF updateCPSR_EnReg = True THEN
                CPSR_Reg_nxt <= flagsFromALU;
            END IF;

            --Handling memory signals if waiting for data from memory to write back to register and wait for memory operation to finish.
            IF writeFromALU_EnReg = False THEN
                procState_nxt <= WRITE_BACK;
                memReadReq    <= '1';
                IF memOpFinished = '1' THEN
                    procState_nxt <= FETCH_SETUP;
                END IF;
            END IF;

            --Handling the actual write backs.
            IF writeBackEnReg = True THEN
                --Load CPSR register.
                IF useCPSR_EnReg = True THEN
                    IF writeFromALU_EnReg = True THEN
                        CPSR_Reg_nxt <= dataFromALU(3 DOWNTO 0);
                    ELSE
                        CPSR_Reg_nxt <= dataFromMem(3 DOWNTO 0);
                    END IF;

                    --Load proper register in register file.
                ELSE
                    loadRegistersSel(destinationRegisterNumberReg) <= '1';
                    IF writeFromALU_EnReg = True THEN
                        dataToRegistersSel <= '0'; --Load registers from ALU output.
                    ELSE
                        dataToRegistersSel <= '1'; --Load register from Memmory.
                    END IF;
                END IF;
            END IF;

            --set ALU signal registers for the next instruction fetch
            operand2SelReg_nxt <= "01111"; --selecting PC as operand 2
            ALU_opCodeReg_nxt  <= "1011";  --tell ALU to MOV PC to output.

        END IF;
    END PROCESS;

    softwareReset <= softwareResetReg;

    --updating registers
    PROCESS (clk, reset)
    BEGIN
        IF reset = '1' THEN
            --control registers
            procState                          <= SETUP;
            instructionReg                     <= (OTHERS => '0');
            CPSR_Reg                           <= (OTHERS => '0');
            CPSR_Reg_Temp                      <= (OTHERS => '0');
            currentlyHandlingInterruptReg      <= False;
            currentlyHandlingInterruptIndexReg <= (OTHERS => '0');
            currentInterruptHandlerAddressReg  <= (OTHERS => '0');
            PC_Reg_Temp                        <= (OTHERS => '0');
            currentlyHaltingReg                <= False;
            invalidInstructionInterruptReg     <= '0';
            softwareInterruptReg               <= '0';

            --registers that to save information about the current instruction
            destinationRegisterNumberReg <= 0;
            addressRegisterNumberReg     <= 0;
            sourceRegisterNumberReg      <= 0;
            useCPSR_EnReg                <= False;
            writeBackEnReg               <= False;
            writeFromALU_EnReg           <= False;
            updateCPSR_EnReg             <= False;
            writeAddressBackEnReg        <= False;
            memOperationReg              <= '0';
            --registers that save the state of the control signals of the ALU
            operand1SelReg           <= (OTHERS => '0');
            operand2SelReg           <= (OTHERS => '0');
            bitManipulationValSelReg <= (OTHERS => '0');
            bitManipulationCodeReg   <= (OTHERS => '0');
            bitManipulationValueReg  <= (OTHERS => '0');

            ALU_opCodeReg <= (OTHERS => '0');
            carryInReg    <= '0';
            upperSelReg   <= '0';
            dataToALU_Reg <= (OTHERS => '0');

            --delay register
            delayReg <= '0';

            softwareResetReg <= '0';

        ELSIF rising_edge(clk) THEN
            IF enable = '1' THEN
                IF alteredClk = '1' THEN
                    --control registers
                    procState                          <= procState_nxt;
                    CPSR_Reg                           <= CPSR_Reg_nxt;
                    CPSR_Reg_Temp                      <= CPSR_Reg_Temp_nxt;
                    PC_Reg_Temp                        <= PC_Reg_Temp_nxt;
                    invalidInstructionInterruptReg     <= invalidInstructionInterruptReg_nxt;
                    softwareInterruptReg               <= softwareInterruptReg_nxt;
                    instructionReg                     <= instructionReg_nxt;
                    currentlyHandlingInterruptReg      <= currentlyHandlingInterruptReg_nxt;
                    currentlyHandlingInterruptIndexReg <= currentlyHandlingInterruptIndexReg_nxt;
                    currentInterruptHandlerAddressReg  <= currentInterruptHandlerAddressReg_nxt;
                    currentlyHaltingReg                <= currentlyHaltingReg_nxt;

                    --registers that to save information about the current instruction
                    destinationRegisterNumberReg <= destinationRegisterNumberReg_nxt;
                    addressRegisterNumberReg     <= addressRegisterNumberReg_nxt;
                    useCPSR_EnReg                <= useCPSR_EnReg_nxt;
                    writeBackEnReg               <= writeBackEnReg_nxt;
                    writeFromALU_EnReg           <= writeFromALU_EnReg_nxt;
                    updateCPSR_EnReg             <= updateCPSR_EnReg_nxt;
                    memOperationReg              <= memOperationReg_nxt;
                    writeAddressBackEnReg        <= writeAddressBackEnReg_nxt;
                    sourceRegisterNumberReg      <= sourceRegisterNumberReg_nxt;

                    --registers that save the state of the control signals of the ALU
                    operand1SelReg           <= operand1SelReg_nxt;
                    operand2SelReg           <= operand2SelReg_nxt;
                    bitManipulationValSelReg <= bitManipulationValSelReg_nxt;
                    bitManipulationCodeReg   <= bitManipulationCodeReg_nxt;
                    bitManipulationValueReg  <= bitManipulationValueReg_nxt;

                    ALU_opCodeReg <= ALU_opCodeReg_nxt;
                    carryInReg    <= carryInReg_nxt;
                    upperSelReg   <= upperSelReg_nxt;
                    dataToALU_Reg <= dataToALU_Reg_nxt;

                    --delay register
                    delayReg <= delayReg_nxt;

                    softwareResetReg <= softwareResetReg_nxt;

                END IF;
            END IF;
        END IF;

    END PROCESS;
END Behavioral;