    signal ram : ram_type :=(
        0 => "11111101",
        1 => "11000000",
        2 => "00000001",
        3 => "01010000",
        4 => "11111101",
        5 => "10000111",
        6 => "11000010",
        7 => "00000000",
        8 => "11111101",
        9 => "10011110",
        10 => "11100000",
        11 => "00000111",
        12 => "11111101",
        13 => "11011111",
        14 => "11111111",
        15 => "11101100",
        others => (others => '0')
    );