    signal ram : ram_type :=(
        0 => "11111101110000000000000101000111",
        others => (others => '0')
    );