    signal ram : ram_type :=(
        0 => "11111101110000000000101000000000",
        1 => "11111101111010000000000000001100",
        2 => "11111001000000000000110000000000",
        3 => "11111101110001001000010010000001",
        4 => "11111101111000000001111010001100",
        5 => "11111001000000000000110000010001",
        6 => "11110000100000000000000000000001",
        7 => "11111101110000000001110101000000",
        8 => "11111101110000000000001000100001",
        9 => "11110000100000000000000000010000",
        10 => "11110000000000000000000000010111",
        11 => "11111011110000000000111101001101",
        12 => "11110110110000000000000000000001",
        13 => "11110100001000000000000000000000",
        14 => "11111101110000000000101010001011",
        15 => "11111101111010000000000000001100",
        16 => "11111001000000000000110010111011",
        17 => "11110000100000000000000010110111",
        18 => "11111101100000000000000110101111",
        others => (others => '0')
    );