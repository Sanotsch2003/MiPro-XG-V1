    signal ram : ram_type :=(
        0 => "11111101110000000000101000001011",
        1 => "11111101111010000000000000001100",
        2 => "11111001000000000000110010111011",
        3 => "11111101110001001000011010001010",
        4 => "11111101111000000001111010001100",
        5 => "11111001000000000000110010101010",
        6 => "11110000100000000000000010111010",
        7 => "11111101110000000000000000000000",
        8 => "11111011110000000000111101001101",
        9 => "11110110110000000000000000101011",
        10 => "11111101110000000000110000001010",
        11 => "11111101111010000000000000001100",
        12 => "11111001000000000000110010101010",
        13 => "11110000000000000000000010101001",
        14 => "11111101100100001000000100101001",
        15 => "11111010111000000000100101000000",
        16 => "00010110011000000000000000000111",
        17 => "11111101110000000000000000000001",
        18 => "11111101110000000000000000000010",
        19 => "11111101110000000000110010001010",
        20 => "11111101111010000000000000001100",
        21 => "11111001000000000000110010101010",
        22 => "11110000000000000000000010101001",
        23 => "11111101110000000010000000001010",
        24 => "11111000001000000000100110100000",
        25 => "00011011110000000000111101001101",
        26 => "00010110110000000000000000010001",
        27 => "11111101110000000001111111101000",
        28 => "11110000100000000000000010101000",
        29 => "11111101110000000000110000001010",
        30 => "11111101111010000000000000001100",
        31 => "11111001000000000000110010101010",
        32 => "11110000000000000000000010101001",
        33 => "11111101100010111000000100101001",
        34 => "00010110011000000000000000000011",
        35 => "11111011010000000000000100110011",
        36 => "11111101100100000110000001100011",
        37 => "11111001000011000110001010010010",
        38 => "11111011110000000000000100010001",
        39 => "11111010111000000000000101000000",
        40 => "00010110011000000000000000010110",
        41 => "11110000100000000000000000000010",
        42 => "11111011110000000000000000010000",
        43 => "11110110011000000000000000100100",
        44 => "11111101110000000000001000001000",
        45 => "11110000100000000000000010101000",
        46 => "11111101110000000000110000001010",
        47 => "11111101111010000000000000001100",
        48 => "11111001000000000000110010101010",
        49 => "11110000000000000000000010101000",
        50 => "11111101100010111000000100001000",
        51 => "00010110011000000000000000000011",
        52 => "11110110011000000000000000101101",
        53 => "11111101110000000000101010000110",
        54 => "11111101111010000000000000001100",
        55 => "11111001000000000000110001100110",
        56 => "11110000100000000000000001100000",
        57 => "11111101100000000000000110101111",
        others => (others => '0')
    );