    signal ram : ram_type :=(
        0 => "11111101110000000000101000001011",
        1 => "11111101111010000000000000001100",
        2 => "11111001000000000000110010111011",
        3 => "11111101110001001000011010001010",
        4 => "11111101111000000001111010001100",
        5 => "11111001000000000000110010101010",
        6 => "11110000100000000000000010111010",
        7 => "11111101110000000000000000000000",
        8 => "11111011110000000000111101001101",
        9 => "11110110110000000000000000011011",
        10 => "11111101110000000000110000001010",
        11 => "11111101111010000000000000001100",
        12 => "11111001000000000000110010101010",
        13 => "11110000000000000000000010101001",
        14 => "11111101100100001000000100101001",
        15 => "11111010111000000000100101000000",
        16 => "00010110011000000000000000000111",
        17 => "11111101110000000000000000000001",
        18 => "11111101110000000000000000000010",
        19 => "11111101110000000000110010001010",
        20 => "11111101111010000000000000001100",
        21 => "11111001000000000000110010101010",
        22 => "11110000000000000000000010101001",
        23 => "11111101110000000010000000001010",
        24 => "11111000001000000000100110100000",
        25 => "00010110010000000000000000010101",
        26 => "11111101100010000110000000100011",
        27 => "11111001000011000110001010010010",
        28 => "11111011110000000000000100010001",
        29 => "11111010111000000000000101000000",
        30 => "00010110011000000000000000001100",
        31 => "11110000100000000000000000000010",
        32 => "11111011110000000000000001000000",
        33 => "11111101110000000001111111101000",
        34 => "11111011110000000000111101001101",
        35 => "11110110110000000000000000000110",
        36 => "11110110011000000000000000011101",
        37 => "11111101110000000000101010000110",
        38 => "11111101111010000000000000001100",
        39 => "11111001000000000000110001100110",
        40 => "11110000100000000000000001100000",
        41 => "11111101100000000000000110101111",
        42 => "11111101110000000000110010000110",
        43 => "11111101111010000000000000001100",
        44 => "11111001000000000000110001100110",
        45 => "11110000100000000000000001101000",
        46 => "11111101100000000000000110101111",
        47 => "11111101110000000001000000001000",
        48 => "11111011110000000000111101001101",
        49 => "11110110111000000000000000001000",
        50 => "11110110011000000000000000101011",
        others => (others => '0')
    );