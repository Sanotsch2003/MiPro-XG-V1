    signal ram : ram_type :=(
        0 => "11111101110000000000110100000000",
        1 => "11111101111010000000000000001100",
        2 => "11111001000000000000110000000000",
        3 => "11111101110000000000001000000001",
        4 => "11110000100000000000000000000001",
        5 => "11111101110000000000110110000000",
        6 => "11111101111010000000000000001100",
        7 => "11111001000000000000110000000000",
        8 => "11111101110000000001111101000001",
        9 => "11110000100000000000000000000001",
        10 => "11111101110000000000111000000000",
        11 => "11111101111010000000000000001100",
        12 => "11111001000000000000110000000000",
        13 => "11111101110000000000000001100001",
        14 => "11110000100000000000000000000001",
        15 => "11111101110000000000111010000000",
        16 => "11111101111010000000000000001100",
        17 => "11111001000000000000110000000000",
        18 => "11111101110000000000010000000001",
        19 => "11110000100000000000000000000001",
        20 => "11111101110000000000111100000000",
        21 => "11111101111010000000000000001100",
        22 => "11111001000000000000110000000000",
        23 => "11111101110111111110000000000001",
        24 => "11110000100000000000000000000001",
        25 => "11111101110000000000111110000000",
        26 => "11111101111010000000000000001100",
        27 => "11111001000000000000110000000000",
        28 => "11111101110000000000000001100001",
        29 => "11110000100000000000000000000001",
        30 => "11111101110000000001000000000000",
        31 => "11111101111010000000000000001100",
        32 => "11111001000000000000110000000000",
        33 => "11111101110000000000100000000001",
        34 => "11110000100000000000000000000001",
        35 => "11111101110000000001000010000000",
        36 => "11111101111010000000000000001100",
        37 => "11111001000000000000110000000000",
        38 => "11111101110101010101010101000001",
        39 => "11110000100000000000000000000001",
        40 => "11111101110000000001000100000000",
        41 => "11111101111010000000000000001100",
        42 => "11111001000000000000110000000000",
        43 => "11111101110000000000000001100001",
        44 => "11110000100000000000000000000001",
        45 => "11111101110000000001000110000000",
        46 => "11111101111010000000000000001100",
        47 => "11111001000000000000110000000000",
        48 => "11111101110000000010000000000001",
        49 => "11110000100000000000000000000001",
        50 => "11111101110000000001001000000000",
        51 => "11111101111010000000000000001100",
        52 => "11111001000000000000110000000000",
        53 => "11111101110000000000000111100001",
        54 => "11110000100000000000000000000001",
        55 => "11111101110000000001001010000000",
        56 => "11111101111010000000000000001100",
        57 => "11111001000000000000110000000000",
        58 => "11111101110000000000000001100001",
        59 => "11110000100000000000000000000001",
        others => (others => '0')
    );