    signal ram : ram_type :=(
        0 => "11111101",
        1 => "11000000",
        2 => "00001010",
        3 => "00000000",
        4 => "11111101",
        5 => "11101000",
        6 => "00000000",
        7 => "00001100",
        8 => "11111001",
        9 => "00000000",
        10 => "00001100",
        11 => "00000000",
        12 => "11111101",
        13 => "11000000",
        14 => "00000000",
        15 => "00000001",
        16 => "11110000",
        17 => "10000000",
        18 => "00000000",
        19 => "00000001",
        20 => "11111101",
        21 => "11000000",
        22 => "00001010",
        23 => "10000000",
        24 => "11111101",
        25 => "11101000",
        26 => "00000000",
        27 => "00001100",
        28 => "11111001",
        29 => "00000000",
        30 => "00001100",
        31 => "00000000",
        32 => "11111101",
        33 => "11000000",
        34 => "00001111",
        35 => "01100001",
        36 => "11110000",
        37 => "10000000",
        38 => "00000000",
        39 => "00000001",
        others => (others => '0')
    );