library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controlUnit is
    Generic(
        numInterrupts : integer := 10
    );

    Port(
        enable                  : in std_logic;
        hardwareReset           : in std_logic;
        softwareReset           : out std_logic;
        clk                     : in std_logic;
        alteredClk              : in std_logic;

        --control signals generated by CU
        operand1Sel             : out std_logic_vector(4 downto 0);
        operand2Sel             : out std_logic_vector(4 downto 0); 
        dataToMemSel            : out std_logic_vector(3 downto 0);

        dataToRegistersSel      : out std_logic;
        loadRegistersSel        : out std_logic_vector(15 downto 0);
        bitManipulationValSel   : out std_logic_vector(4 downto 0);

        bitManipulationCode     : out std_logic_vector(1 downto 0);
        bitManipulationValue    : out std_logic_vector(4 downto 0);

        ALU_opCode              : out std_logic_vector(3 downto 0);
        carryIn                 : out std_logic;
        upperSel                : out std_logic;

        memWriteReq             : out std_logic;
        memReadReq              : out std_logic;

        clearInterrupts         : out std_logic_vector(numInterrupts-1 downto 0);
        dataToALU               : out std_logic_vector(31 downto 0);

        ALU_En                  : out std_logic;
          
        --signals controlling the CU
        programmingMode         : in std_logic;
        IVT_address             : in std_logic_vector(31 downto 0);
        dataFromMem             : in std_logic_vector(31 downto 0);
        dataFromALU             : in std_logic_vector(31 downto 0);
        flagsFromALU            : in std_logic_vector(3 downto 0);
        memOpFinished           : in std_logic;
        --debug signals
        debug : out std_logic_vector(49 downto 0)
);
end controlUnit;

architecture Behavioral of controlUnit is
    --type StateType      is (SETUP, FETCH1, FETCH2, FETCH3, FETCH4, DECODE, EXECUTE, MEMORY_ACCESS, WRITE_BACK);

    --signal state        : StateType    := FETCH1;
    --signal state_nxt    : StateType;
    
    type procStateType is (SETUP, FETCH_SETUP, FETCH_MEM_READ, DECODE, EXECUTE, MEM_ACCESS, WRITE_BACK);
    --type executeStateType is (DECODE_EXECUTE1, DECODE_EXECUTE2);
    
    signal procState, procState_nxt : procStateType;
    --signal executeState, executeState_nxt : executeStateType;


    --internal registers
    signal currentlyHandlingInterruptReg, currentlyHandlingInterruptReg_nxt : boolean;
    signal currentlyHaltingReg, currentlyHaltingReg_nxt : boolean;

    signal softwareResetReg, softwareResetReg_nxt : std_logic;

    --signals to keep track of decoded information within instructions
    signal instructionReg, instructionReg_nxt : std_logic_vector(31 downto 0);
    signal destinationRegisterNumberReg, destinationRegisterNumberReg_nxt : integer;
    signal addressRegisterNumberReg, addressRegisterNumberReg_nxt : integer;
    signal sourceRegisterNumberReg, sourceRegisterNumberReg_nxt : integer;
    signal useCPSR_EnReg, useCPSR_EnReg_nxt : boolean;
    signal writeBackEnReg, writeBackEnReg_nxt : boolean;
    signal writeFromALU_EnReg, writeFromALU_EnReg_nxt : boolean;
    signal updateCPSR_EnReg, updateCPSR_EnReg_nxt : boolean;
    signal writeAddressBackEnReg, writeAddressBackEnReg_nxt : boolean;
    signal memOperationReg, memOperationReg_nxt : std_logic; --1: read, 0: write

    signal CPSR_Reg                      : std_logic_vector(3 downto 0);
    signal CPSR_Reg_nxt                  : std_logic_vector(3 downto 0);

    signal Z_flag : std_logic;
    signal N_flag : std_logic;
    signal V_flag : std_logic;
    signal C_flag : std_logic; 

    --registers that keep track of the control signals of the ALU (only the control Signal for the ALU need a separate register) 
    signal operand1SelReg, operand1SelReg_nxt                       : std_logic_vector(4 downto 0) := (others => '0');
    signal operand2SelReg, operand2SelReg_nxt                       : std_logic_vector(4 downto 0) := (others => '0');
    signal bitManipulationValSelReg, bitManipulationValSelReg_nxt   : std_logic_vector(4 downto 0) := (others => '0');
    signal bitManipulationCodeReg, bitManipulationCodeReg_nxt       : std_logic_vector(1 downto 0) := (others => '0');
    signal bitManipulationValueReg, bitManipulationValueReg_nxt     : std_logic_vector(4 downto 0) := (others => '0');

    signal ALU_opCodeReg, ALU_opCodeReg_nxt                         : std_logic_vector(3 downto 0) := (others => '0');
    signal carryInReg, carryInReg_nxt                               : std_logic := '0';
    signal upperSelReg, upperSelReg_nxt                             : std_logic := '0';
    signal dataToALU_Reg, dataToALU_Reg_nxt                           : std_logic_vector(31 downto 0) := (others => '0');

    --delay register
    signal delayReg, delayReg_nxt : std_logic;

    --interrupt register
    signal invalidInstructionInterruptReg, invalidInstructionInterruptReg_nxt   : std_logic;
    signal softwareInterruptReg, softwareInterruptReg_nxt : std_logic;

    --Shift register for detecting rising edge of the programming mode signal.
    signal programmingModeShiftReg : std_logic_vector(1 downto 0);


    --bit masks
    type bitMasksType is array (0 to 16) of std_logic_vector(31 downto 0);

    constant bitMasks : bitMasksType :=(
        0 => x"00000000",
        1 => x"00000001",
        2 => x"00000003",
        3 => x"0000000F",
        4 => x"000000FF",
        5 => x"0000FF00",
        6 => x"0F0F0F0F",
        7 => x"F0F0F0F0",
        8 => x"55555555",
        9 => x"AAAAAAAA",
        10 => x"FFFFFFFF",
        others => (others => '0')
    );

    --operation codes
    --Data Processing
    constant ANDD: std_logic_vector(3 downto 0) := "0000";
    constant EOR: std_logic_vector(3 downto 0) := "0001";
    constant ORR: std_logic_vector(3 downto 0) := "0010";
    constant BIC: std_logic_vector(3 downto 0) := "0011";
    constant NOTT: std_logic_vector(3 downto 0) := "0100";
    constant SUB: std_logic_vector(3 downto 0) := "0101";
    constant BUSS: std_logic_vector(3 downto 0) := "0110";
    constant ADDD: std_logic_vector(3 downto 0) := "0111";
    constant ADC: std_logic_vector(3 downto 0) := "1000";
    constant SBC: std_logic_vector(3 downto 0) := "1001";
    constant BSC: std_logic_vector(3 downto 0) := "1010";
    constant MOV: std_logic_vector(3 downto 0) := "1011";
    constant MUL: std_logic_vector(3 downto 0) := "1100";
    constant UMUL: std_logic_vector(3 downto 0) := "1101";

    --Data Movement 
    constant LOAD : std_logic_vector(2 downto 0) := "000";
    constant STORE: std_logic_vector(2 downto 0) := "001";

    --Special Instructions
    constant PASS : std_logic_vector(3 downto 0) := "0000";
    constant HALT: std_logic_vector(3 downto 0) := "0001";
    constant SIR : std_logic_vector(3 downto 0) := "0010";
    constant RES : std_logic_vector(3 downto 0) := "0011";


    --Control Flow 

    --Booloader code. This code is executed when programming mode is enabled.
    type ROM is array (0 to 256) of std_logic_vector(31 downto 0);
    signal bootloaderMemory : ROM :=(
        0 => "11111101110000000000101000001011",
        1 => "11111101111010000000000000001100",
        2 => "11111001000000000000110010111011",
        3 => "11111101110001001000011010001010",
        4 => "11111101111000000001111010001100",
        5 => "11111001000000000000110010101010",
        6 => "11110000100000000000000010111010",
        7 => "11111101110000000000000000000000",
        8 => "11111011110000000000111101001101",
        9 => "11110110110000000000000000011011",
        10 => "11111101110000000000110000001010",
        11 => "11111101111010000000000000001100",
        12 => "11111001000000000000110010101010",
        13 => "11110000000000000000000010101001",
        14 => "11111101100100001000000100101001",
        15 => "11111010111000000000100101000000",
        16 => "00010110011000000000000000000111",
        17 => "11111101110000000000000000000001",
        18 => "11111101110000000000000000000010",
        19 => "11111101110000000000110010001010",
        20 => "11111101111010000000000000001100",
        21 => "11111001000000000000110010101010",
        22 => "11110000000000000000000010101001",
        23 => "11111101110000000010000000001010",
        24 => "11111000001000000000100110100000",
        25 => "00010110010000000000000000010101",
        26 => "11111101100010000110000000100011",
        27 => "11111001000011000110001010010010",
        28 => "11111011110000000000000100010001",
        29 => "11111010111000000000000101000000",
        30 => "00010110011000000000000000001100",
        31 => "11110000100000000000000000000010",
        32 => "11111011110000000000000001000000",
        33 => "11111101110000000001111111101000",
        34 => "11111011110000000000111101001101",
        35 => "11110110110000000000000000000110",
        36 => "11110110011000000000000000011101",
        37 => "11111101110000000000101010000110",
        38 => "11111101111010000000000000001100",
        39 => "11111001000000000000110001100110",
        40 => "11110000100000000000000001100000",
        41 => "11111101100000000000000110101111",
        42 => "11111101110000000000110010000110",
        43 => "11111101111010000000000000001100",
        44 => "11111001000000000000110001100110",
        45 => "11110000100000000000000001101000",
        46 => "11111101100000000000000110101111",
        47 => "11111101110000000001000000001000",
        48 => "11111011110000000000111101001101",
        49 => "11110110111000000000000000001000",
        50 => "11110110011000000000000000101011",
        others => (others => '0')
    );
    
begin
    Z_flag <= CPSR_Reg(3);
    N_flag <= CPSR_Reg(2);
    V_flag <= CPSR_Reg(1);
    C_flag <= CPSR_Reg(0);

    softwareReset <= softwareResetReg;

    stateMachine : process(procState, operand1SelReg, operand2SelReg, bitManipulationValSelReg, bitManipulationCodeReg, bitManipulationValueReg, ALU_opCodeReg, carryInReg, upperSelReg, dataToALU_Reg, programmingMode, IVT_address, dataFromMem, dataFromALU, flagsFromALU, memOpFinished, instructionReg, destinationRegisterNumberReg, useCPSR_EnReg, writeBackEnReg, writeFromALU_EnReg, updateCPSR_EnReg, memOperationReg, addressRegisterNumberReg, writeAddressBackEnReg, sourceRegisterNumberReg, CPSR_Reg, Z_flag, N_flag, V_flag, C_flag, softwareInterruptReg, invalidInstructionInterruptReg, currentlyHandlingInterruptReg, currentlyHaltingReg, delayReg, softwareResetReg)
        variable condition          : std_logic_vector(3 downto 0);
        variable conditionMet       : std_logic;
        type instructionClassType is (DATA_PROCESSING, DATA_MOVEMENT, SPECIAL, CONTROL_FLOW, INVALID); 
        variable instructionClass : instructionClassType;

        --variables for the different instruction classes:
        --Data Processing
        variable dataProcessingOpCode : std_logic_vector(3 downto 0);

        --Data Movement
        variable dataMovementOpCode : std_logic_vector(2 downto 0);

        --Special Instructions
        variable specialInstructionOpCode : std_logic_vector(3 downto 0);

        --Control Flow
        variable controlFlowOpCode : std_logic_vector(1 downto 0);

        --variables for different sections within the instruction:
        variable sourceReg      : std_logic_vector(3 downto 0);
        variable addressRegister: std_logic_vector(3 downto 0);
        variable immediateEn    : std_logic;
        variable offsetEn       : std_logic;
        variable offset         : std_logic_vector(11 downto 0);
        variable subtractEn     : std_logic;
        variable immediateValue : std_logic_vector(31 downto 0);

        variable bitManipulationMethod : std_logic_vector(1 downto 0);
        variable bitManipulationUseRegEn : std_logic;
        variable bitManipulationOperand : std_logic_vector(4 downto 0);
        
    begin
        --default assignments for control signals
        operand1Sel                         <= (others => '1');
        operand2Sel                         <= (others => '1');
        dataToMemSel                        <= (others => '0');
        dataToRegistersSel                  <= '0';
        bitManipulationValSel               <= (others => '1');
        loadRegistersSel                    <= (others => '0');
        bitManipulationCode                 <= (others => '0');
        bitManipulationValue                <= (others => '0');
        ALU_opCode                          <= (others => '0');
        carryIn                             <= '0';
        upperSel                            <= '0';
        memWriteReq                         <= '0';
        memReadReq                          <= '0';
        clearInterrupts                     <= (others => '0');
        dataToALU                           <= (others => '0');
        ALU_En                              <= '0';

        --controlRegisters
        instructionReg_nxt                  <= instructionReg;
        procState_nxt                       <= procState;
        CPSR_Reg_nxt                        <= CPSR_Reg;
        invalidInstructionInterruptReg_nxt  <= invalidInstructionInterruptReg;
        softwareInterruptReg_nxt            <= softwareInterruptReg;
        currentlyHandlingInterruptReg_nxt   <= currentlyHandlingInterruptReg;
        currentlyHaltingReg_nxt             <= currentlyHaltingReg;

        --temporary registers for holding information about the current instruction
        destinationRegisterNumberReg_nxt    <= destinationRegisterNumberReg;
        addressRegisterNumberReg_nxt        <= addressRegisterNumberReg;
        useCPSR_EnReg_nxt                   <= useCPSR_EnReg;
        writeBackEnReg_nxt                  <= writeBackEnReg;
        writeFromALU_EnReg_nxt              <= writeFromALU_EnReg;
        updateCPSR_EnReg_nxt                <= updateCPSR_EnReg; 
        memOperationReg_nxt                 <= memOperationReg;
        writeAddressBackEnReg_nxt           <= writeAddressBackEnReg;
        sourceRegisterNumberReg_nxt         <= sourceRegisterNumberReg;

        --registers that save the state of the control signals of the ALU
        operand1SelReg_nxt                  <= operand1SelReg;
        operand2SelReg_nxt                  <= operand2SelReg;
        bitManipulationValSelReg_nxt        <= bitManipulationValSelReg;
        bitManipulationCodeReg_nxt          <= bitManipulationCodeReg;
        bitManipulationValueReg_nxt         <= bitManipulationValueReg;
        ALU_opCodeReg_nxt                   <= ALU_opCodeReg;
        carryInReg_nxt                      <= carryInReg;
        upperSelReg_nxt                     <= upperSelReg;
        dataToALU_Reg_nxt                   <= dataToALU_Reg;  
        
        --delay register
        delayReg_nxt                        <= delayReg;

        --reset register
        softwareResetReg_nxt                <= softwareResetReg;
        
        if procState = SETUP then
            procState_nxt       <= FETCH_SETUP;
            --set ALU signal registers for the next instruction fetch
            operand2SelReg_nxt         <= "01111";     --selecting PC as operand 2
            ALU_opCodeReg_nxt          <= "1011";      --tell ALU to MOV PC to output.

        elsif procState = FETCH_SETUP then
            if currentlyHaltingReg = False then
                procState_nxt       <= FETCH_MEM_READ;

                --set ALU control signals
                operand2Sel         <= operand2SelReg;
                ALU_opCode          <= ALU_opCodeReg;  

                --enable ALU
                ALU_En              <= '1'; 

                --Prepare ALU control signals for next state, where the PC will be incremented.
                operand1SelReg_nxt         <= "10000";                 --dataToALU as operand 1.
                operand2SelReg_nxt         <= "01111";                 --Selecting PC as operand 2.
                dataToALU_Reg_nxt           <= x"00000004";             --set dataToALU to 4 to increment PC later
                ALU_opCodeReg_nxt          <= "0111";                  --tell ALU to add operand1 (4) to the PC
            else
                procState_nxt <= FETCH_SETUP;
            end if;

        elsif procState = FETCH_MEM_READ then
            memReadReq          <= '1';
            operand1Sel         <= operand1SelReg;
            operand2Sel         <= operand2SelReg;
            dataToALU           <= dataToALU_Reg;
            ALU_opCode          <= ALU_opCodeReg;
            --Handle instruction fetch in programming mode.
            if programmingMode = '1' then
                instructionReg_nxt  <= bootloaderMemory(to_integer(unsigned(dataFromALU(9 downto 2)))); --Address needs to be divided by four.
                ALU_En <= '1';                              --enable ALU in order to increment the PC
                procState_nxt <= DECODE;

            --Handle instruction fetch in normal mode.
            else
                if memOpFinished = '1' then                     --wait for data to arrive         
                    instructionReg_nxt  <= dataFromMem;         --load current instruction into the instruction register
                    ALU_En <= '1';                              --enable ALU in order to increment the PC
                    procState_nxt <= DECODE;
                end if;
            end if;


        elsif procState = DECODE then
            --this instruction is also used to write the updated instruction address back to the PC
            loadRegistersSel    <= "1000000000000000";  --load value back into PC
            dataToRegistersSel  <= '0';         --sending data from ALU to registers in order to write the incremented address back to the PC

            procState_nxt <= EXECUTE; --The next state will always be "EXECUTE" state.

            --default assignments
            operand1SelReg_nxt                  <= (others => '0');
            operand2SelReg_nxt                  <= (others => '0');
            bitManipulationValSelReg_nxt        <= (others => '1');
            bitManipulationCodeReg_nxt          <= (others => '0');
            bitManipulationValueReg_nxt         <= (others => '0');
            ALU_opCodeReg_nxt                   <= (others => '0');
            carryInReg_nxt                      <= '0'; --not used yet
            upperSelReg_nxt                     <= '0'; --not used yet
            dataToALU_Reg_nxt                    <= (others => '0');     

            --extract condition from instruction
            condition := instructionReg(31 downto 28);
            case condition is
                when "0000" => conditionMet := Z_flag;                                  --equal
                when "0001" => conditionMet := not Z_flag;                              --not equal
                when "0010" => conditionMet := C_flag;                                  --unsigned higher or same
                when "0011" => conditionMet := not C_flag;                              --unsigned lower
                when "0100" => conditionMet := N_flag;                                  --negative
                when "0101" => conditionMet := not N_flag;                              --positive or zero
                when "0110" => conditionMet := V_flag;                                  --overflow
                when "1101" => conditionMet := (not Z_flag) or (N_flag xor V_flag);     --less than or equal
                when others => conditionMet := '1';                                     --always
            end case;
            
            --skip instruction if condition is not met
            if not conditionMet = '1' then
                --set ALU signal registers for the next instruction fetch
                operand2SelReg_nxt         <= "01111";     --selecting PC as operand 2
                ALU_opCodeReg_nxt          <= "1011";      --tell ALU to MOV PC to output.
                procState_nxt <= FETCH_SETUP; 
            else
                --IF an instruction uses bit manipulation, it will ALWAYS use bit 20-13. Therefore, it can be set in the beginning without any conditions. However, each instruction sets "bitManipulationValSel" individually depending on whether (and if yes how) it  uses bit manipulation. Setting "bitManipulationValSel="11111"" will tell the ALU to not make use of bit manipulation.
                bitManipulationMethod            := instructionReg(20 downto 19);
                bitManipulationUseRegEn          := instructionReg(18);
                bitManipulationOperand           := instructionReg(17 downto 13);
                bitManipulationCodeReg_nxt       <= bitManipulationMethod;
                bitManipulationValueReg_nxt      <= bitManipulationOperand;

                --check what kind of instruction class the instruction belongs to
                if instructionReg(27) = '1' then
                    instructionClass := DATA_PROCESSING;
                elsif instructionReg(27 downto 26) = "00" then
                    instructionClass := DATA_MOVEMENT;
                elsif instructionReg(27 downto 25) = "010" then
                    instructionClass := SPECIAL;
                elsif instructionReg(27 downto 25) = "011" then
                    instructionClass := CONTROL_FLOW;
                else
                    instructionClass := INVALID; --needs to be set to avoid latch
                    invalidInstructionInterruptReg_nxt <= '1'; --handle invalid instructions
                    procState_nxt <= SETUP;
                end if;

            
                --handle different instructin classes 
                case instructionClass is
                    when DATA_PROCESSING =>
                        updateCPSR_EnReg_nxt <= True;--All of the Data Processing instructions update the CPSR register.
                        useCPSR_EnReg_nxt <= False; --this is a default assignments, in some cases the CPSR will be used as the destination register.
                        writeBackEnReg_nxt <= True; --This instruction class always writes back to register file.
                        writeFromALU_EnReg_nxt <= True; --This instruction class updates registers from ALU result.

                        destinationRegisterNumberReg_nxt <= to_integer(unsigned(instructionReg(3 downto 0))); --All instructions in this instruction class use the same bits for the destination Register.
                        
                        immediateEn := instructionReg(22);--All instructions in this instruction class use the same bit as their "Immediate Enable Bit".
                        
                        dataProcessingOpCode := instructionReg(26 downto 23);
                        ALU_opCodeReg_nxt <= dataProcessingOpCode; --Tell ALU which operation to perform.
                        
                        if dataProcessingOpCode = MOV then --the MOV instruction is different from the other ones.
                            if instructionReg(4) = '1' then --if this bit is set, the destination register is the CPSR.
                                useCPSR_EnReg_nxt <= True;
                            end if;
                            
                            if immediateEn = '1' then 
                                if instructionReg(21) = '1' then --checks if the "Load Higher Bytes Enable Bit" is set.
                                    immediateValue := instructionReg(20 downto 5) & x"0000";
                                else
                                    immediateValue := x"0000" & instructionReg(20 downto 5);
                                end if;
                                operand2SelReg_nxt <= "10000"; --tells the ALU to use "dataToALU" as operand 2.
                                dataToALU_Reg_nxt <= immediateValue;
                            else
                                operand2SelReg_nxt <= instructionReg(9 downto 5);
                                if instructionReg(9) = '1' then --if this bit is set, the source register is the CPSR.
                                    dataToALU_Reg_nxt <= x"0000000" & CPSR_Reg;
                                end if;
                                if bitManipulationUseRegEn = '0' then 
                                    bitManipulationValSelReg_nxt <= "10000"; --uses the "bitManipulationOperand" as immediate value for bit manipulation.
                                else
                                    bitManipulationValSelReg_nxt <= '0' & bitManipulationOperand(3 downto 0); --uses the "bitManipulationOperand" as register for bit manipulation
                                end if;
                            
                            end if;
                        else
                            --all of these instruction will always apply bit manipulation to operand 2
                            if bitManipulationUseRegEn = '0' then 
                                bitManipulationValSelReg_nxt <= "10000"; --uses the "bitManipulationOperand" as immediate value for bit manipulation.
                            else
                                bitManipulationValSelReg_nxt <= '0' & bitManipulationOperand(3 downto 0); --uses the "bitManipulationOperand" as register for bit manipulation
                            end if;
    
                            --all instruction specify the operand 1 register in the same way
                            operand1SelReg_nxt <= '0' & instructionReg(11 downto 8);
    
                            --all instructions use the same bit to tell the cpu, if operand 2 should be interpreted as a register or as something else.      
                            if immediateEn = '1' then
                                operand2SelReg_nxt <= "10000"; --operand 2 will be specified by CU
                            else 
                                operand2SelReg_nxt <= '0' & instructionReg(7 downto 4); --operand 2 will be a register
                            end if;
    
    
                            if dataProcessingOpCode = ANDD or dataProcessingOpCode = EOR or dataProcessingOpCode = ORR or dataProcessingOpCode = BIC or dataProcessingOpCode = NOTT then
                                --These instructions do not offer the possibility to specify immediate values. Instead, a bit mask can be specified.
                                if immediateEn = '1' then
                                    dataToALU_Reg_nxt <= bitMasks(to_integer(unsigned(instructionReg(7 downto 4))));
                                end if;
                                --These instructions can disable write back if bit 21 of the instruction is set.
                                if instructionReg(21) = '1' then
                                    writeBackEnReg_nxt <= False;
                                end if;

                            elsif dataProcessingOpCode = SUB or dataProcessingOpCode = BUSS or dataProcessingOpCode = ADDD or dataProcessingOpCode = ADC or dataProcessingOpCode = SBC or dataProcessingOpCode = BSC then
                                --These instructions offer you to specify an immediate value.
                                if immediateEn = '1' then
                                    dataToALU_Reg_nxt <= x"0000000" & instructionReg(7 downto 4);
                                end if;

                                --These instructions can disable write back if bit 21 of the instruction is set.
                                if instructionReg(21) = '1' then
                                    writeBackEnReg_nxt <= False;
                                end if;

                            elsif dataProcessingOpCode = MUL or dataProcessingOpCode = UMUL then 
                                --These instructions offer you to specify an immediate value.
                                if immediateEn = '1' then
                                    dataToALU_Reg_nxt <= x"0000000" & instructionReg(7 downto 4);
                                end if;
                                --Since these instructions perform multiplications, it needs to be specified, whether to write back the upper or lower 32 bits of the result.
                                upperSelReg_nxt <= instructionReg(21);
                            else
                                invalidInstructionInterruptReg_nxt <= '1';
                            end if;

                        end if;
                        
                    
                    when DATA_MOVEMENT =>
                        dataMovementOpCode := instructionReg(25 downto 23);
                        updateCPSR_EnReg_nxt <= False;--None of the Data Processing instructions update the CPSR register.
                        useCPSR_EnReg_nxt <= False; --None of the Data Movement instructions update the status flags.
                        writeBackEnReg_nxt <= True; --This instruction class always updates the registers.
                        writeFromALU_EnReg_nxt <= False; --This instruction class updates registers from memory.
                        writeAddressBackEnReg_nxt <= False; --This is a default assignment. In some cases the altered address will be written back to the addressRegister.

                        if dataMovementOpCode = STORE or dataMovementOpCode = LOAD then
                            --differentiate between load and store instruction
                            if dataMovementOpCode = STORE then
                                memOperationReg_nxt <= '0';
                                sourceRegisterNumberReg_nxt <= to_integer(unsigned(instructionReg(3 downto 0))); --CAN BE REMOVED???
                            else
                                memOperationReg_nxt <= '1';
                                destinationRegisterNumberReg_nxt <= to_integer(unsigned(instructionReg(3 downto 0)));
                            end if;

                            --otherwise, the two instructions work exactly the same:
                            addressRegister := instructionReg(7 downto 4);
                            addressRegisterNumberReg_nxt <= to_integer(unsigned(addressRegister));
                            operand2SelReg_nxt <= '0' & addressRegister; --operand 2 will be data in specified register.
                            operand1SelReg_nxt <= "10000"; --operand one will be the data sent by control unit.

                            offsetEn := instructionReg(21);
                            if offsetEn = '1' then
                                subtractEn := instructionReg(20);
                                offset     := instructionReg(19 downto 8);
                                dataToALU_Reg_nxt  <= x"00000" & offset;
                                --subtract or add the offset to the current
                                if subtractEn = '1' then
                                    ALU_opCodeReg_nxt <= "0110"; --operation code for subraction (operand2 - operand1)
                                else
                                    ALU_opCodeReg_nxt <= "0111"; --operation code for addition (operand2 + operand 1)
                                end if;
                            else
                                --ignore operand 1
                                ALU_opCodeReg_nxt <= "1011";
                                --Apply bit manipulation to operand2.
                                if bitManipulationUseRegEn = '0' then 
                                    bitManipulationValSelReg_nxt <= "10000"; --Uses the "bitManipulationOperand" as immediate value for bit manipulation.
                                else
                                    bitManipulationValSelReg_nxt <= '0' & bitManipulationOperand(3 downto 0); --uses the "bitManipulationOperand" as register for bit manipulation.
                                end if;   
                            end if;
                            if instructionReg(22) = '1' then
                                writeAddressBackEnReg_nxt <= True;
                            end if;
                        else
                            invalidInstructionInterruptReg_nxt <= '1'; --handle invalid instructions
                            procState_nxt <= SETUP; 
                        end if;
                    
                    when SPECIAL =>
                        specialInstructionOpCode := instructionReg(24 downto 21);
                        updateCPSR_EnReg_nxt <= False;--None of the Data Processing instructions update the CPSR register.
                        useCPSR_EnReg_nxt <= False; --None of the Data Movement instructions update the status flags.
                        writeBackEnReg_nxt <= False; --This instruction class never updates the registers.
                        
                        --None of these instruction need memory access and they do not write back to the register file.
                        --Set ALU signal registers for the next instruction fetch.
                        operand2SelReg_nxt         <= "01111";     --Selecting PC as operand 2
                        ALU_opCodeReg_nxt          <= "1011";      --Tell ALU to MOV PC to output.
                        --Go to next instruction
                        procState_nxt <= FETCH_SETUP; 

                        case specialInstructionOpCode is 
                        when PASS =>
                            null;
                        when HALT =>
                            currentlyHaltingReg_nxt <= True;

                        when SIR =>
                            softwareInterruptReg_nxt <= '1';
                        when RES =>
                            softwareResetReg_nxt <= '1';
                        when others =>
                            invalidInstructionInterruptReg_nxt <= '1'; --Handle invalid instructions.
                            procState_nxt <= SETUP;
                        end case;

                    when CONTROL_FLOW =>
                        controlFlowOpCode := instructionReg(24 downto 23);
                        updateCPSR_EnReg_nxt <= False;--None of the Data Processing instructions update the CPSR register.
                        useCPSR_EnReg_nxt <= False; --None of the Data Movement instructions update the status flags.
                        writeBackEnReg_nxt <= True; --This instruction class always updates the registers.
                        writeFromALU_EnReg_nxt <= True; --This instruction class updates registers from the ALU.
                                   
                        --The program counter is always the source register 
                        destinationRegisterNumberReg_nxt <= 15;

                        --set the ALU signals
                        operand1SelReg_nxt <= "01111"; --Select PC as operand 1.
                        if instructionReg(22) = '1' then --Check if 'Immediate Offset Enable Bit' is set.
                            operand2SelReg_nxt <= "10000"; --Select data from CU as operand 2.
                            dataToALU_Reg_nxt <= "000000000" & instructionReg(20 downto 0) & "00";  --Multiply immediate value by 4 (so that it is a valid memory address) and send it to ALU.
                            if instructionReg(21) = '1' then --Check if the 'Subtract Bit' is set.
                                ALU_opCodeReg_nxt <= "0101"; --ALU operation Code for subtraction.
                            else
                                ALU_opCodeReg_nxt <= "0111"; --ALU operation Code for addition.
                            end if;
                        else
                            operand2SelReg_nxt <= '0' & instructionReg(3 downto 0); --Select specified register as operand 2.
                            if bitManipulationUseRegEn = '0' then 
                                bitManipulationValSelReg_nxt <= "10000"; --uses the "bitManipulationOperand" as immediate value for bit manipulation.
                            else
                                bitManipulationValSelReg_nxt <= '0' & bitManipulationOperand(3 downto 0); --uses the "bitManipulationOperand" as register for bit manipulation
                            end if;
                            if instructionReg(21) = '1' then --Check if the 'Register as Offset Enable Bit' is set.
                                ALU_opCodeReg_nxt <= "0111"; --ALU operation Code for addition (offset will be added to the PC)
                            else
                                ALU_opCodeReg_nxt <= "1011"; --ALU operation Code for MOV (The value of operand2 will be copied into the PC).
                            end if;
                        end if;
                        
                    when others =>
                        invalidInstructionInterruptReg_nxt <= '1'; --Handle invalid instructions.
                        procState_nxt <= SETUP;
                end case;
            end if;

        elsif procState = Execute then
            ALU_En                  <= '1'; --enable ALU
            operand1Sel             <= operand1SelReg;
            operand2Sel             <= operand2SelReg;
            bitManipulationValSel   <= bitManipulationValSelReg;
            bitManipulationCode     <= bitManipulationCodeReg;
            bitManipulationValue    <= bitManipulationValueReg;
            ALU_opCode              <= ALU_opCodeReg;
            carryIn                 <= carryInReg;
            upperSel                <= upperSelReg;
            dataToALU               <= dataToALU_Reg;

            --wait one clock cycle for the result and the flags to arrive
            if delayReg = '1' then
                if writeFromALU_EnReg = True then
                    procState_nxt <= WRITE_BACK;
                else
                    procState_nxt <= MEM_ACCESS;
                end if;
                delayReg_nxt <= '0';
            else
                delayReg_nxt <= '1';
            end if;

        
        elsif procState = MEM_ACCESS then
            if memOperationReg = '1' then --read
                memReadReq <= '1';
                procState_nxt <= WRITE_BACK; --After loading a value from memory, that value needs to be written to a register. 
            else
                memWriteReq <= '1'; --write
                if memOpFinished = '1' then
                    procState_nxt <= FETCH_SETUP; --After storing a value in memory, No register access will be needed.
                end if;
            end if;
            dataToMemSel <= std_logic_vector(to_unsigned(sourceRegisterNumberReg, 4)); 
            
            if writeAddressBackEnReg = True then 
                loadRegistersSel(addressRegisterNumberReg) <= '1'; --Select address register as write back register.
                dataToRegistersSel <= '0'; --Load registers from ALU output.
            end if;

            --set ALU signal registers for the next instruction fetch
            operand2SelReg_nxt         <= "01111";     --selecting PC as operand 2
            ALU_opCodeReg_nxt          <= "1011";      --tell ALU to MOV PC to output.
            
        elsif procState = WRITE_BACK then
            --default assignment
            procState_nxt <= FETCH_SETUP;

            --Handling the updates of the status flags.
            if updateCPSR_EnReg = True then
                CPSR_Reg_nxt <= flagsFromALU; 
            end if;

            --Handling memory signals if waiting for data from memory to write back to register and wait for memory operation to finish.
            if writeFromALU_EnReg = False then
                procState_nxt <= WRITE_BACK;
                memReadReq <= '1';
                if memOpFinished = '1' then
                    procState_nxt <= FETCH_SETUP;
                end if;
            end if;

            --Handling the actual write backs.
            if writeBackEnReg = True then
                --Load CPSR register.
                if useCPSR_EnReg = True then
                    if writeFromALU_EnReg = True then
                        CPSR_Reg_nxt <= dataFromALU(3 downto 0); 
                    else
                        CPSR_Reg_nxt <= dataFromMem(3 downto 0);
                    end if;
                    
                 --Load proper register in register file.
                else
                    loadRegistersSel(destinationRegisterNumberReg) <= '1';
                    if writeFromALU_EnReg = True then
                        dataToRegistersSel <= '0'; --Load registers from ALU output.
                    else
                        dataToRegistersSel <= '1'; --Load register from Memmory.
                    end if;
                end if;
       

            end if;

            --set ALU signal registers for the next instruction fetch
            operand2SelReg_nxt         <= "01111";     --selecting PC as operand 2
            ALU_opCodeReg_nxt          <= "1011";      --tell ALU to MOV PC to output.

        end if;
    end process;


    --updating registers
    process(clk, hardwareReset, softwareResetReg)
        variable programmingModeShiftRegVariable : std_logic_vector(1 downto 0);
    begin
        if hardwareReset = '1' or softwareResetReg = '1' then
            --control registers
            procState                       <= SETUP;
            instructionReg                  <= (others => '0');
            CPSR_Reg                        <= (others => '0');
            currentlyHandlingInterruptReg   <= False;
            currentlyHaltingReg             <= False;
            invalidInstructionInterruptReg  <= '0';
            softwareInterruptReg            <= '0';

            --registers that to save information about the current instruction
            destinationRegisterNumberReg <= 0;
            addressRegisterNumberReg <= 0;
            sourceRegisterNumberReg <= 0;
            useCPSR_EnReg <= False;
            writeBackEnReg <= False;
            writeFromALU_EnReg <= False;
            updateCPSR_EnReg <= False;
            writeAddressBackEnReg <= False;
            memOperationReg <= '0';


            --registers that save the state of the control signals of the ALU
            operand1SelReg                  <= (others => '0');
            operand2SelReg                  <= (others => '0');
            bitManipulationValSelReg        <= (others => '0');
            bitManipulationCodeReg          <= (others => '0');
            bitManipulationValueReg         <= (others => '0');

            ALU_opCodeReg                   <= (others => '0');
            carryInReg                      <= '0';
            upperSelReg                     <= '0';
            dataToALU_Reg                   <= (others => '0');

            --delay register
            delayReg                        <= '0';

            --reset register                
            softwareResetReg                <= '0';
            
            if hardwareReset = '1' then 
                programmingModeShiftReg <= "00";
            end if;

            
        elsif rising_edge(clk) then
            if enable = '1' then
                if alteredClk = '1' then
                    --control registers
                    procState                       <= procState_nxt;
                    CPSR_Reg                        <= CPSR_Reg_nxt;
                    invalidInstructionInterruptReg  <= invalidInstructionInterruptReg_nxt;
                    softwareInterruptReg            <= softwareInterruptReg_nxt;
                    instructionReg                  <= instructionReg_nxt;
                    currentlyHandlingInterruptReg   <= currentlyHandlingInterruptReg_nxt;
                    currentlyHaltingReg             <= currentlyHaltingReg_nxt;

                    --registers that to save information about the current instruction
                    destinationRegisterNumberReg    <= destinationRegisterNumberReg_nxt;
                    addressRegisterNumberReg        <= addressRegisterNumberReg_nxt;
                    useCPSR_EnReg                   <= useCPSR_EnReg_nxt;
                    writeBackEnReg                  <= writeBackEnReg_nxt;
                    writeFromALU_EnReg              <= writeFromALU_EnReg_nxt;
                    updateCPSR_EnReg                <= updateCPSR_EnReg_nxt; 
                    memOperationReg                 <= memOperationReg_nxt;
                    writeAddressBackEnReg           <= writeAddressBackEnReg_nxt;
                    sourceRegisterNumberReg         <= sourceRegisterNumberReg_nxt;

                    --registers that save the state of the control signals of the ALU
                    operand1SelReg                  <= operand1SelReg_nxt;
                    operand2SelReg                  <= operand2SelReg_nxt;
                    bitManipulationValSelReg        <= bitManipulationValSelReg_nxt;
                    bitManipulationCodeReg          <= bitManipulationCodeReg_nxt;
                    bitManipulationValueReg         <= bitManipulationValueReg_nxt;

                    ALU_opCodeReg                   <= ALU_opCodeReg_nxt;
                    carryInReg                      <= carryInReg_nxt;
                    upperSelReg                     <= upperSelReg_nxt;
                    dataToALU_Reg                   <= dataToALU_Reg_nxt;      

                    --delay register
                    delayReg                        <= delayReg_nxt;

                    --reset register
                    softwareResetReg                <= softwareResetReg_nxt;
                    
                    --Shift register for detecting rising edge of debug mode signal
                    programmingModeShiftRegVariable := programmingModeShiftReg(0) & programmingMode;
                    programmingModeShiftReg <= programmingModeShiftRegVariable;
                    --Reset processor on rising and falling edge of programming mode signal.
                    if programmingModeShiftRegVariable = "01" or programmingModeShiftRegVariable = "10" then
                        softwareResetReg <= '1';
                    end if;
                    
                end if;
            end if;
        end if;

    end process;


end Behavioral;
