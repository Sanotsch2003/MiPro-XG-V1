this is a tet
