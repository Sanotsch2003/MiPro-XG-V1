library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity RAM is
    generic(
        ramSize : integer
    );
    port (
        enable                     : in std_logic;
        clk                        : in std_logic;
        reset                      : in std_logic;
        alteredClk                 : in std_logic;
        address                    : in std_logic_vector(31 downto 0);
        dataIn                     : in std_logic_vector(31 downto 0);
        dataOut                    : out std_logic_vector(31 downto 0);
        writeEn                    : in std_logic;
        readEn                     : in std_logic;
        memOpFinished              : out std_logic
    );
end RAM;

architecture Behavioral of RAM is
    type ram_type is array (0 to ramSize-1) of std_logic_vector(31 downto 0);
    
    --deafult count program
    signal ram : ram_type :=(
        0 => "11111101110000000001010110000000",
        1 => "11111101111010000000000000001100",
        2 => "11111001000000000000110000000000",
        3 => "11111101110000000000000000100001",
        4 => "11110000100000000000000000000001",
        5 => "11111101110000000001011110000000",
        6 => "11111101111010000000000000001100",
        7 => "11111001000000000000110000000000",
        8 => "11111101110000000000000000100001",
        9 => "11110000100000000000000000000001",
        10 => "11111101110000000001100110000000",
        11 => "11111101111010000000000000001100",
        12 => "11111001000000000000110000000000",
        13 => "11111101110000000000000000100001",
        14 => "11110000100000000000000000000001",
        15 => "11111101110000000001101110000000",
        16 => "11111101111010000000000000001100",
        17 => "11111001000000000000110000000000",
        18 => "11111101110000000000000000000001",
        19 => "11110000100000000000000000000001",
        20 => "11111101110000000001110110000000",
        21 => "11111101111010000000000000001100",
        22 => "11111001000000000000110000000000",
        23 => "11111101110000000000000000000001",
        24 => "11110000100000000000000000000001",
        25 => "11111101110000000001111110000000",
        26 => "11111101111010000000000000001100",
        27 => "11111001000000000000110000000000",
        28 => "11111101110000000000000000000001",
        29 => "11110000100000000000000000000001",
        30 => "11111101110000000010000110000000",
        31 => "11111101111010000000000000001100",
        32 => "11111001000000000000110000000000",
        33 => "11111101110000000000000000000001",
        34 => "11110000100000000000000000000001",
        35 => "11111101110000000010001110000000",
        36 => "11111101111010000000000000001100",
        37 => "11111001000000000000110000000000",
        38 => "11111101110000000000000000000001",
        39 => "11110000100000000000000000000001",
        40 => "11111101110000000010010110000000",
        41 => "11111101111010000000000000001100",
        42 => "11111001000000000000110000000000",
        43 => "11111101110000000000000000000001",
        44 => "11110000100000000000000000000001",
        45 => "11111101110000000010011110000000",
        46 => "11111101111010000000000000001100",
        47 => "11111001000000000000110000000000",
        48 => "11111101110000000000000000000001",
        49 => "11110000100000000000000000000001",
        50 => "11111101110000000010100110000000",
        51 => "11111101111010000000000000001100",
        52 => "11111001000000000000110000000000",
        53 => "11111101110000000000000000000001",
        54 => "11110000100000000000000000000001",
        55 => "11111101110000000010101110000000",
        56 => "11111101111010000000000000001100",
        57 => "11111001000000000000110000000000",
        58 => "11111101110000000000000000000001",
        59 => "11110000100000000000000000000001",
        60 => "11111101110000000010110110000000",
        61 => "11111101111010000000000000001100",
        62 => "11111001000000000000110000000000",
        63 => "11111101110000000000000000000001",
        64 => "11110000100000000000000000000001",
        65 => "11111101110000000010111110000000",
        66 => "11111101111010000000000000001100",
        67 => "11111001000000000000110000000000",
        68 => "11111101110000000000000000000001",
        69 => "11110000100000000000000000000001",
        70 => "11111101110000000011000110000000",
        71 => "11111101111010000000000000001100",
        72 => "11111001000000000000110000000000",
        73 => "11111101110000000000000000000001",
        74 => "11110000100000000000000000000001",
        75 => "11111101110000000011001110000000",
        76 => "11111101111010000000000000001100",
        77 => "11111001000000000000110000000000",
        78 => "11111101110000000000000000000001",
        79 => "11110000100000000000000000000001",
        others => (others => '0')
    );
  
begin
    process(clk, reset) 
    begin 
        if rising_edge(clk) then 
            --if alteredClk = '1' then
                if writeEn = '1' then
                    -- Write data to RAM
                    ram(to_integer(unsigned(address))) <= dataIn;
                end if;
        
                if readEn = '1' then
                    -- Read data from RAM
                    dataOut <= ram(to_integer(unsigned(address)));
                else
                    dataOut <= (others => '0');
                    
                end if;
            --end if;
        end if;

    end process;
    
    --Setting the memOpFinished signal.
    process(clk)
    begin
        if rising_edge(clk) then
            --if alteredClk = '1' then
                if writeEn = '1' or readEn = '1' then
                    memOpFinished <= '1';
                else
                    memOpFinished <= '0';
                end if;
            --end if;
        end if;
    end process;

end Behavioral;
