    signal ram : ram_type :=(
        0 => "11111101110000000000101000000000",
        1 => "11111101111010000000000000001100",
        2 => "11111001000000000000110000000000",
        3 => "11111101110001001000010010000111",
        4 => "11111101111000000001111010001100",
        5 => "11111001000000000000110001110111",
        6 => "11110000110000000000000000000111",
        7 => "11111101110000000000101010000000",
        8 => "11111101111010000000000000001100",
        9 => "11111001000000000000110000000000",
        10 => "11111101110000101100010111000111",
        11 => "11110000110000000000000000000111",
        12 => "11110100001000000000000000000000",
        others => (others => '0')
    );