    signal ram : ram_type :=(
        0 => "11111011110000000000111101001101",
        1 => "11110110110000000000000000000101",
        2 => "11111101110000001001101001001011",
        3 => "11111101110000000000000001100000",
        4 => "11111011110000000000111101001101",
        5 => "11110110110000000000000000000001",
        6 => "11110110011000000000000000000100",
        7 => "11111101110000000000000001100001",
        8 => "11111010101000000000000100000000",
        9 => "00001101100000000000000110101111",
        others => (others => '0')
    );